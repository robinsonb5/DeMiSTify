library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8ecc287",
    12 => x"48c0c44e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90588",
    17 => x"49d8ecc2",
    18 => x"48e4d7c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"e4d7c287",
    25 => x"e0d7c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e1c187f7",
    29 => x"d7c287c1",
    30 => x"d7c24de4",
    31 => x"ad744ce4",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"c04b710e",
    37 => x"9a4a134c",
    38 => x"7287cd02",
    39 => x"87e0c049",
    40 => x"4a1384c1",
    41 => x"87f3059a",
    42 => x"4c264874",
    43 => x"4f264b26",
    44 => x"8148731e",
    45 => x"c502a973",
    46 => x"05531287",
    47 => x"4f2687f6",
    48 => x"c0ff1e1e",
    49 => x"c4486a4a",
    50 => x"a6c498c0",
    51 => x"02987058",
    52 => x"7a7187f3",
    53 => x"4f262648",
    54 => x"ff1e731e",
    55 => x"ffc34bd4",
    56 => x"c34a6b7b",
    57 => x"496b7bff",
    58 => x"b17232c8",
    59 => x"6b7bffc3",
    60 => x"7131c84a",
    61 => x"7bffc3b2",
    62 => x"32c8496b",
    63 => x"4871b172",
    64 => x"4d2687c4",
    65 => x"4b264c26",
    66 => x"5e0e4f26",
    67 => x"0e5d5c5b",
    68 => x"d4ff4a71",
    69 => x"c348724c",
    70 => x"7c7098ff",
    71 => x"bfe4d7c2",
    72 => x"d087c805",
    73 => x"30c94866",
    74 => x"d058a6d4",
    75 => x"29d84966",
    76 => x"ffc34871",
    77 => x"d07c7098",
    78 => x"29d04966",
    79 => x"ffc34871",
    80 => x"d07c7098",
    81 => x"29c84966",
    82 => x"ffc34871",
    83 => x"d07c7098",
    84 => x"ffc34866",
    85 => x"727c7098",
    86 => x"7129d049",
    87 => x"98ffc348",
    88 => x"4b6c7c70",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87fffd",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487dffd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c1fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87defc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"49e3c878",
   125 => x"d387d5fa",
   126 => x"c01ec04b",
   127 => x"c1c1f0ff",
   128 => x"87c6fc49",
   129 => x"987086c4",
   130 => x"ff87ca05",
   131 => x"ffc348d4",
   132 => x"cb48c178",
   133 => x"87ebfd87",
   134 => x"ff058bc1",
   135 => x"48c087db",
   136 => x"4387e3fb",
   137 => x"5300444d",
   138 => x"20434844",
   139 => x"6c696166",
   140 => x"49000a21",
   141 => x"00525245",
   142 => x"00495053",
   143 => x"74697257",
   144 => x"61662065",
   145 => x"64656c69",
   146 => x"5e0e000a",
   147 => x"ff0e5c5b",
   148 => x"eefc4cd4",
   149 => x"1eeac687",
   150 => x"c1f0e1c0",
   151 => x"e9fa49c8",
   152 => x"c186c487",
   153 => x"87c802a8",
   154 => x"c087fdfd",
   155 => x"87e8c148",
   156 => x"7087e5f9",
   157 => x"ffffcf49",
   158 => x"a9eac699",
   159 => x"fd87c802",
   160 => x"48c087e6",
   161 => x"c387d1c1",
   162 => x"f1c07cff",
   163 => x"87c7fc4b",
   164 => x"c0029870",
   165 => x"1ec087eb",
   166 => x"c1f0ffc0",
   167 => x"e9f949fa",
   168 => x"7086c487",
   169 => x"87d90598",
   170 => x"6c7cffc3",
   171 => x"7cffc349",
   172 => x"c17c7c7c",
   173 => x"c40299c0",
   174 => x"db48c187",
   175 => x"d748c087",
   176 => x"05abc287",
   177 => x"e7c887ca",
   178 => x"87c0f749",
   179 => x"87c848c0",
   180 => x"fe058bc1",
   181 => x"48c087f7",
   182 => x"0e87e9f8",
   183 => x"5d5c5b5e",
   184 => x"d0ff1e0e",
   185 => x"c0c0c84d",
   186 => x"e4d7c24b",
   187 => x"c878c148",
   188 => x"d7f649f8",
   189 => x"6d4cc787",
   190 => x"c4987348",
   191 => x"987058a6",
   192 => x"6d87cc02",
   193 => x"c4987348",
   194 => x"987058a6",
   195 => x"c287f405",
   196 => x"87eff97d",
   197 => x"9873486d",
   198 => x"7058a6c4",
   199 => x"87cc0298",
   200 => x"9873486d",
   201 => x"7058a6c4",
   202 => x"87f40598",
   203 => x"1ec07dc3",
   204 => x"c1d0e5c0",
   205 => x"d1f749c0",
   206 => x"c186c487",
   207 => x"87c105a8",
   208 => x"05acc24c",
   209 => x"f3c887cb",
   210 => x"87c0f549",
   211 => x"cec148c0",
   212 => x"058cc187",
   213 => x"fb87e0fe",
   214 => x"d7c287f0",
   215 => x"987058e8",
   216 => x"c187cd05",
   217 => x"f0ffc01e",
   218 => x"f649d0c1",
   219 => x"86c487dc",
   220 => x"c348d4ff",
   221 => x"ddc578ff",
   222 => x"ecd7c287",
   223 => x"73486d58",
   224 => x"58a6c498",
   225 => x"cc029870",
   226 => x"73486d87",
   227 => x"58a6c498",
   228 => x"f4059870",
   229 => x"ff7dc287",
   230 => x"ffc348d4",
   231 => x"2648c178",
   232 => x"0e87dff5",
   233 => x"5d5c5b5e",
   234 => x"c0c81e0e",
   235 => x"4cc04bc0",
   236 => x"dfcdeec5",
   237 => x"5ca6c44a",
   238 => x"c34cd4ff",
   239 => x"486c7cff",
   240 => x"05a8fec3",
   241 => x"7187c0c2",
   242 => x"e2c00599",
   243 => x"bfd0ff87",
   244 => x"c4987348",
   245 => x"987058a6",
   246 => x"ff87ce02",
   247 => x"7348bfd0",
   248 => x"58a6c498",
   249 => x"f2059870",
   250 => x"48d0ff87",
   251 => x"d478d1c4",
   252 => x"b7c04866",
   253 => x"e0c006a8",
   254 => x"7cffc387",
   255 => x"99714a6c",
   256 => x"7187c702",
   257 => x"0a7a970a",
   258 => x"66d481c1",
   259 => x"d888c148",
   260 => x"b7c058a6",
   261 => x"e0ff01a8",
   262 => x"7cffc387",
   263 => x"0599717c",
   264 => x"ff87e1c0",
   265 => x"7348bfd0",
   266 => x"58a6c498",
   267 => x"ce029870",
   268 => x"bfd0ff87",
   269 => x"c4987348",
   270 => x"987058a6",
   271 => x"ff87f205",
   272 => x"78d048d0",
   273 => x"c17e4ac1",
   274 => x"eefd058a",
   275 => x"26486e87",
   276 => x"0e87eff2",
   277 => x"0e5c5b5e",
   278 => x"c84a711e",
   279 => x"c04bc0c0",
   280 => x"48d4ff4c",
   281 => x"ff78ffc3",
   282 => x"7348bfd0",
   283 => x"58a6c498",
   284 => x"ce029870",
   285 => x"bfd0ff87",
   286 => x"c4987348",
   287 => x"987058a6",
   288 => x"ff87f205",
   289 => x"c3c448d0",
   290 => x"48d4ff78",
   291 => x"7278ffc3",
   292 => x"f0ffc01e",
   293 => x"f149d1c1",
   294 => x"86c487f0",
   295 => x"c0059870",
   296 => x"c0c887ee",
   297 => x"4966d41e",
   298 => x"c487f8fb",
   299 => x"ff4c7086",
   300 => x"7348bfd0",
   301 => x"58a6c498",
   302 => x"ce029870",
   303 => x"bfd0ff87",
   304 => x"c4987348",
   305 => x"987058a6",
   306 => x"ff87f205",
   307 => x"78c248d0",
   308 => x"f0264874",
   309 => x"5e0e87ee",
   310 => x"0e5d5c5b",
   311 => x"ffc01ec0",
   312 => x"49c9c1f0",
   313 => x"d287e3f0",
   314 => x"f2d7c21e",
   315 => x"87f3fa49",
   316 => x"4cc086c8",
   317 => x"b7d284c1",
   318 => x"87f804ac",
   319 => x"97f2d7c2",
   320 => x"c0c349bf",
   321 => x"a9c0c199",
   322 => x"87e7c005",
   323 => x"97f9d7c2",
   324 => x"31d049bf",
   325 => x"97fad7c2",
   326 => x"32c84abf",
   327 => x"d7c2b172",
   328 => x"4abf97fb",
   329 => x"cf4c71b1",
   330 => x"9cffffff",
   331 => x"34ca84c1",
   332 => x"c287e7c1",
   333 => x"bf97fbd7",
   334 => x"c631c149",
   335 => x"fcd7c299",
   336 => x"c74abf97",
   337 => x"b1722ab7",
   338 => x"97f7d7c2",
   339 => x"cf4d4abf",
   340 => x"f8d7c29d",
   341 => x"c34abf97",
   342 => x"c232ca9a",
   343 => x"bf97f9d7",
   344 => x"7333c24b",
   345 => x"fad7c2b2",
   346 => x"c34bbf97",
   347 => x"b7c69bc0",
   348 => x"c2b2732b",
   349 => x"7148c181",
   350 => x"c1497030",
   351 => x"70307548",
   352 => x"c14c724d",
   353 => x"c8947184",
   354 => x"06adb7c0",
   355 => x"34c187cc",
   356 => x"c0c82db7",
   357 => x"ff01adb7",
   358 => x"487487f4",
   359 => x"0e87e3ed",
   360 => x"0e5c5b5e",
   361 => x"4cc04b71",
   362 => x"c04866d0",
   363 => x"c006a8b7",
   364 => x"4a1387e3",
   365 => x"bf9766cc",
   366 => x"4866cc49",
   367 => x"a6d080c1",
   368 => x"aab77158",
   369 => x"c187c402",
   370 => x"c187cc48",
   371 => x"b766d084",
   372 => x"ddff04ac",
   373 => x"c248c087",
   374 => x"264d2687",
   375 => x"264b264c",
   376 => x"5b5e0e4f",
   377 => x"c20e5d5c",
   378 => x"c048d8e0",
   379 => x"d0d8c278",
   380 => x"f949c01e",
   381 => x"86c487dd",
   382 => x"c5059870",
   383 => x"c848c087",
   384 => x"4bc087ef",
   385 => x"48d0e5c2",
   386 => x"1ec878c1",
   387 => x"1efde0c0",
   388 => x"49c6d9c2",
   389 => x"c887c8fe",
   390 => x"05987086",
   391 => x"e5c287c6",
   392 => x"78c048d0",
   393 => x"e1c01ec8",
   394 => x"d9c21ec6",
   395 => x"eefd49e2",
   396 => x"7086c887",
   397 => x"87c60598",
   398 => x"48d0e5c2",
   399 => x"e5c278c0",
   400 => x"c002bfd0",
   401 => x"dfc287fa",
   402 => x"c24bbfd6",
   403 => x"bf9fcee0",
   404 => x"ead6c54a",
   405 => x"87c705aa",
   406 => x"bfd6dfc2",
   407 => x"ca87cc4b",
   408 => x"02aad5e9",
   409 => x"48c087c5",
   410 => x"c287c6c7",
   411 => x"731ed0d8",
   412 => x"87dff749",
   413 => x"987086c4",
   414 => x"c087c505",
   415 => x"87f1c648",
   416 => x"e1c01ec8",
   417 => x"d9c21ecf",
   418 => x"d2fc49e2",
   419 => x"7086c887",
   420 => x"87c80598",
   421 => x"48d8e0c2",
   422 => x"87da78c1",
   423 => x"e1c01ec8",
   424 => x"d9c21ed8",
   425 => x"f6fb49c6",
   426 => x"7086c887",
   427 => x"c5c00298",
   428 => x"c548c087",
   429 => x"e0c287fb",
   430 => x"49bf97ce",
   431 => x"05a9d5c1",
   432 => x"c287cdc0",
   433 => x"bf97cfe0",
   434 => x"a9eac249",
   435 => x"87c5c002",
   436 => x"dcc548c0",
   437 => x"d0d8c287",
   438 => x"c34cbf97",
   439 => x"c002ace9",
   440 => x"ebc387cc",
   441 => x"c5c002ac",
   442 => x"c548c087",
   443 => x"d8c287c3",
   444 => x"49bf97db",
   445 => x"ccc00599",
   446 => x"dcd8c287",
   447 => x"c249bf97",
   448 => x"c5c002a9",
   449 => x"c448c087",
   450 => x"d8c287e7",
   451 => x"48bf97dd",
   452 => x"58d4e0c2",
   453 => x"e0c288c1",
   454 => x"d8c258d8",
   455 => x"49bf97de",
   456 => x"d8c28173",
   457 => x"4abf97df",
   458 => x"7135c84d",
   459 => x"f0e4c285",
   460 => x"e0d8c25d",
   461 => x"c248bf97",
   462 => x"c258c4e5",
   463 => x"02bfd8e0",
   464 => x"c887dcc2",
   465 => x"f4e0c01e",
   466 => x"e2d9c21e",
   467 => x"87cff949",
   468 => x"987086c8",
   469 => x"87c5c002",
   470 => x"d4c348c0",
   471 => x"d0e0c287",
   472 => x"c4484abf",
   473 => x"e0e0c230",
   474 => x"c0e5c258",
   475 => x"f5d8c25a",
   476 => x"c849bf97",
   477 => x"f4d8c231",
   478 => x"a14bbf97",
   479 => x"f6d8c249",
   480 => x"d04bbf97",
   481 => x"49a17333",
   482 => x"97f7d8c2",
   483 => x"33d84bbf",
   484 => x"c249a173",
   485 => x"c259c8e5",
   486 => x"91bfc0e5",
   487 => x"bfece4c2",
   488 => x"f4e4c281",
   489 => x"fdd8c259",
   490 => x"c84bbf97",
   491 => x"fcd8c233",
   492 => x"a34cbf97",
   493 => x"fed8c24b",
   494 => x"d04cbf97",
   495 => x"4ba37434",
   496 => x"97ffd8c2",
   497 => x"9ccf4cbf",
   498 => x"a37434d8",
   499 => x"f8e4c24b",
   500 => x"738bc25b",
   501 => x"f8e4c292",
   502 => x"78a17248",
   503 => x"c287cbc1",
   504 => x"bf97e2d8",
   505 => x"c231c849",
   506 => x"bf97e1d8",
   507 => x"c249a14a",
   508 => x"c559e0e0",
   509 => x"81ffc731",
   510 => x"e5c229c9",
   511 => x"d8c259c0",
   512 => x"4abf97e7",
   513 => x"d8c232c8",
   514 => x"4bbf97e6",
   515 => x"e5c24aa2",
   516 => x"e5c25ac8",
   517 => x"7592bfc0",
   518 => x"fce4c282",
   519 => x"f4e4c25a",
   520 => x"c278c048",
   521 => x"7248f0e4",
   522 => x"49c078a1",
   523 => x"c187f7c7",
   524 => x"87e5f648",
   525 => x"33544146",
   526 => x"20202032",
   527 => x"54414600",
   528 => x"20203631",
   529 => x"41460020",
   530 => x"20323354",
   531 => x"46002020",
   532 => x"32335441",
   533 => x"00202020",
   534 => x"31544146",
   535 => x"20202036",
   536 => x"5b5e0e00",
   537 => x"710e5d5c",
   538 => x"d8e0c24a",
   539 => x"87cc02bf",
   540 => x"b7c74b72",
   541 => x"c14d722b",
   542 => x"87ca9dff",
   543 => x"b7c84b72",
   544 => x"c34d722b",
   545 => x"d8c29dff",
   546 => x"e4c21ed0",
   547 => x"7349bfec",
   548 => x"feee7181",
   549 => x"7086c487",
   550 => x"87c50598",
   551 => x"e6c048c0",
   552 => x"d8e0c287",
   553 => x"87d202bf",
   554 => x"91c44975",
   555 => x"81d0d8c2",
   556 => x"ffcf4c69",
   557 => x"9cffffff",
   558 => x"497587cb",
   559 => x"d8c291c2",
   560 => x"699f81d0",
   561 => x"f448744c",
   562 => x"5e0e87cf",
   563 => x"0e5d5c5b",
   564 => x"4c7186f4",
   565 => x"e5c24bc0",
   566 => x"c47ebfc8",
   567 => x"e5c248a6",
   568 => x"c878bfcc",
   569 => x"78c048a6",
   570 => x"bfdce0c2",
   571 => x"06a8c048",
   572 => x"c887ddc2",
   573 => x"99cf4966",
   574 => x"c287d805",
   575 => x"c81ed0d8",
   576 => x"c1484966",
   577 => x"58a6cc80",
   578 => x"c487c8ed",
   579 => x"d0d8c286",
   580 => x"c087c34b",
   581 => x"6b9783e0",
   582 => x"c1029a4a",
   583 => x"e5c387e1",
   584 => x"dac102aa",
   585 => x"49a3cb87",
   586 => x"d8496997",
   587 => x"cec10599",
   588 => x"c01ecb87",
   589 => x"731e66e0",
   590 => x"87e3f149",
   591 => x"987086c8",
   592 => x"87fbc005",
   593 => x"c44aa3dc",
   594 => x"796a49a4",
   595 => x"c849a3da",
   596 => x"699f4da4",
   597 => x"e0c27d48",
   598 => x"d302bfd8",
   599 => x"49a3d487",
   600 => x"c049699f",
   601 => x"7199ffff",
   602 => x"c430d048",
   603 => x"87c258a6",
   604 => x"486e7ec0",
   605 => x"7d70806d",
   606 => x"48c17cc0",
   607 => x"c887c5c1",
   608 => x"80c14866",
   609 => x"c258a6cc",
   610 => x"a8bfdce0",
   611 => x"87e3fd04",
   612 => x"bfd8e0c2",
   613 => x"87eac002",
   614 => x"c4fb496e",
   615 => x"58a6c487",
   616 => x"ffcf4970",
   617 => x"99f8ffff",
   618 => x"87d602a9",
   619 => x"89c24970",
   620 => x"bfd0e0c2",
   621 => x"f0e4c291",
   622 => x"807148bf",
   623 => x"fc58a6c8",
   624 => x"48c087e1",
   625 => x"d0f08ef4",
   626 => x"1e731e87",
   627 => x"496a4a71",
   628 => x"7a7181c1",
   629 => x"bfd4e0c2",
   630 => x"87cb0599",
   631 => x"6b4ba2c8",
   632 => x"87fdf949",
   633 => x"c17b4970",
   634 => x"87f1ef48",
   635 => x"711e731e",
   636 => x"f0e4c24b",
   637 => x"a3c849bf",
   638 => x"c24a6a4a",
   639 => x"d0e0c28a",
   640 => x"a17292bf",
   641 => x"d4e0c249",
   642 => x"9a6b4abf",
   643 => x"c849a172",
   644 => x"e8711e66",
   645 => x"86c487fd",
   646 => x"c4059870",
   647 => x"c248c087",
   648 => x"ee48c187",
   649 => x"5e0e87f7",
   650 => x"710e5c5b",
   651 => x"724bc04a",
   652 => x"e0c0029a",
   653 => x"49a2da87",
   654 => x"c24b699f",
   655 => x"02bfd8e0",
   656 => x"a2d487cf",
   657 => x"49699f49",
   658 => x"ffffc04c",
   659 => x"c234d09c",
   660 => x"744cc087",
   661 => x"029b73b3",
   662 => x"c24a87df",
   663 => x"d0e0c28a",
   664 => x"c29249bf",
   665 => x"48bff0e4",
   666 => x"e5c28072",
   667 => x"487158d0",
   668 => x"e0c230c4",
   669 => x"e9c058e0",
   670 => x"f4e4c287",
   671 => x"e5c24bbf",
   672 => x"e4c248cc",
   673 => x"c278bff8",
   674 => x"02bfd8e0",
   675 => x"e0c287c9",
   676 => x"c449bfd0",
   677 => x"c287c731",
   678 => x"49bffce4",
   679 => x"e0c231c4",
   680 => x"e5c259e0",
   681 => x"f2ec5bcc",
   682 => x"5b5e0e87",
   683 => x"f40e5d5c",
   684 => x"9a4a7186",
   685 => x"c287de02",
   686 => x"c048ccd8",
   687 => x"c4d8c278",
   688 => x"cce5c248",
   689 => x"d8c278bf",
   690 => x"e5c248c8",
   691 => x"c078bfc8",
   692 => x"c048fff1",
   693 => x"dce0c278",
   694 => x"d8c249bf",
   695 => x"714abfcc",
   696 => x"cbc403aa",
   697 => x"cf497287",
   698 => x"e0c00599",
   699 => x"d0d8c287",
   700 => x"c4d8c21e",
   701 => x"d8c249bf",
   702 => x"a1c148c4",
   703 => x"d2e57178",
   704 => x"c086c487",
   705 => x"c248fbf1",
   706 => x"cc78d0d8",
   707 => x"fbf1c087",
   708 => x"e0c048bf",
   709 => x"fff1c080",
   710 => x"ccd8c258",
   711 => x"80c148bf",
   712 => x"58d0d8c2",
   713 => x"000c7b27",
   714 => x"bf97bf00",
   715 => x"c2029c4c",
   716 => x"e5c387ee",
   717 => x"e7c202ac",
   718 => x"fbf1c087",
   719 => x"a3cb4bbf",
   720 => x"cf4d1149",
   721 => x"d6c105ad",
   722 => x"df497487",
   723 => x"cd89c199",
   724 => x"e0e0c291",
   725 => x"4aa3c181",
   726 => x"a3c35112",
   727 => x"c551124a",
   728 => x"51124aa3",
   729 => x"124aa3c7",
   730 => x"4aa3c951",
   731 => x"a3ce5112",
   732 => x"d051124a",
   733 => x"51124aa3",
   734 => x"124aa3d2",
   735 => x"4aa3d451",
   736 => x"a3d65112",
   737 => x"d851124a",
   738 => x"51124aa3",
   739 => x"124aa3dc",
   740 => x"4aa3de51",
   741 => x"f1c05112",
   742 => x"78c148ff",
   743 => x"7587c1c1",
   744 => x"0599c849",
   745 => x"7587f3c0",
   746 => x"0599d049",
   747 => x"66dc87d0",
   748 => x"87cac002",
   749 => x"66dc4973",
   750 => x"0298700f",
   751 => x"f1c087dc",
   752 => x"c005bfff",
   753 => x"e0c287c6",
   754 => x"50c048e0",
   755 => x"48fff1c0",
   756 => x"f1c078c0",
   757 => x"c248bffb",
   758 => x"f1c087dc",
   759 => x"78c048ff",
   760 => x"bfdce0c2",
   761 => x"ccd8c249",
   762 => x"aa714abf",
   763 => x"87f5fb04",
   764 => x"bfcce5c2",
   765 => x"87c8c005",
   766 => x"bfd8e0c2",
   767 => x"87f4c102",
   768 => x"bfc8d8c2",
   769 => x"87d9f149",
   770 => x"58ccd8c2",
   771 => x"e0c27e70",
   772 => x"c002bfd8",
   773 => x"496e87dd",
   774 => x"ffffffcf",
   775 => x"02a999f8",
   776 => x"c487c8c0",
   777 => x"78c048a6",
   778 => x"c487e6c0",
   779 => x"78c148a6",
   780 => x"6e87dec0",
   781 => x"f8ffcf49",
   782 => x"c002a999",
   783 => x"a6c887c8",
   784 => x"c078c048",
   785 => x"a6c887c5",
   786 => x"c478c148",
   787 => x"66c848a6",
   788 => x"0566c478",
   789 => x"6e87ddc0",
   790 => x"c289c249",
   791 => x"91bfd0e0",
   792 => x"bff0e4c2",
   793 => x"c2807148",
   794 => x"c258c8d8",
   795 => x"c048ccd8",
   796 => x"87e1f978",
   797 => x"8ef448c0",
   798 => x"0087dee5",
   799 => x"00000000",
   800 => x"1e000000",
   801 => x"c348d4ff",
   802 => x"496878ff",
   803 => x"87c60299",
   804 => x"05a9fbc0",
   805 => x"487187ee",
   806 => x"5e0e4f26",
   807 => x"710e5c5b",
   808 => x"ff4bc04a",
   809 => x"ffc348d4",
   810 => x"99496878",
   811 => x"87c1c102",
   812 => x"02a9ecc0",
   813 => x"c087fac0",
   814 => x"c002a9fb",
   815 => x"66cc87f3",
   816 => x"cc03abb7",
   817 => x"0266d087",
   818 => x"097287c7",
   819 => x"c1097997",
   820 => x"02997182",
   821 => x"83c187c2",
   822 => x"c348d4ff",
   823 => x"496878ff",
   824 => x"87cd0299",
   825 => x"02a9ecc0",
   826 => x"fbc087c7",
   827 => x"cdff05a9",
   828 => x"0266d087",
   829 => x"97c087c3",
   830 => x"a9fbc07a",
   831 => x"7387c705",
   832 => x"8c0cc04c",
   833 => x"4c7387c2",
   834 => x"87c24874",
   835 => x"4c264d26",
   836 => x"4f264b26",
   837 => x"48d4ff1e",
   838 => x"6878ffc3",
   839 => x"b7f0c049",
   840 => x"87ca04a9",
   841 => x"a9b7f9c0",
   842 => x"c087c301",
   843 => x"c1c189f0",
   844 => x"ca04a9b7",
   845 => x"b7c6c187",
   846 => x"87c301a9",
   847 => x"7189f7c0",
   848 => x"0e4f2648",
   849 => x"5d5c5b5e",
   850 => x"7186f40e",
   851 => x"4bd4ff4c",
   852 => x"c37e4dc0",
   853 => x"d0ff7bff",
   854 => x"c0c848bf",
   855 => x"a6c898c0",
   856 => x"02987058",
   857 => x"d0ff87d0",
   858 => x"c0c848bf",
   859 => x"a6c898c0",
   860 => x"05987058",
   861 => x"d0ff87f0",
   862 => x"78e1c048",
   863 => x"c2fc7bd4",
   864 => x"99497087",
   865 => x"87c7c102",
   866 => x"c87bffc3",
   867 => x"786b48a6",
   868 => x"c04866c8",
   869 => x"c802a8fb",
   870 => x"e8e5c287",
   871 => x"eec002bf",
   872 => x"714dc187",
   873 => x"e6c00299",
   874 => x"a9fbc087",
   875 => x"fb87c302",
   876 => x"ffc387d1",
   877 => x"c1496b7b",
   878 => x"cc05a9c6",
   879 => x"7bffc387",
   880 => x"48a6c87b",
   881 => x"49c0786b",
   882 => x"0599714d",
   883 => x"7587daff",
   884 => x"dec1059d",
   885 => x"7bffc387",
   886 => x"ffc34a6b",
   887 => x"48a6c47b",
   888 => x"486e786b",
   889 => x"a6c480c1",
   890 => x"49a4c858",
   891 => x"c8496997",
   892 => x"da05a966",
   893 => x"49a4c987",
   894 => x"aa496997",
   895 => x"ca87d005",
   896 => x"699749a4",
   897 => x"a966c449",
   898 => x"c187c405",
   899 => x"c887d64d",
   900 => x"ecc04866",
   901 => x"87c902a8",
   902 => x"c04866c8",
   903 => x"c405a8fb",
   904 => x"c17ec087",
   905 => x"7bffc34d",
   906 => x"6b48a6c8",
   907 => x"029d7578",
   908 => x"ff87e2fe",
   909 => x"c848bfd0",
   910 => x"c898c0c0",
   911 => x"987058a6",
   912 => x"ff87d002",
   913 => x"c848bfd0",
   914 => x"c898c0c0",
   915 => x"987058a6",
   916 => x"ff87f005",
   917 => x"e0c048d0",
   918 => x"f4486e78",
   919 => x"87ecfa8e",
   920 => x"5c5b5e0e",
   921 => x"86f40e5d",
   922 => x"ff59a6c4",
   923 => x"c0c84cd0",
   924 => x"1e6e4bc0",
   925 => x"49ece5c2",
   926 => x"c487cfe9",
   927 => x"02987086",
   928 => x"c287f7c5",
   929 => x"4dbff0e5",
   930 => x"f6fa496e",
   931 => x"58a6c887",
   932 => x"9873486c",
   933 => x"7058a6cc",
   934 => x"87cc0298",
   935 => x"9873486c",
   936 => x"7058a6c4",
   937 => x"87f40598",
   938 => x"d4ff7cc5",
   939 => x"78d5c148",
   940 => x"bfe8e5c2",
   941 => x"c481c149",
   942 => x"8ac14a66",
   943 => x"487232c6",
   944 => x"d4ffb071",
   945 => x"486c7808",
   946 => x"a6c49873",
   947 => x"02987058",
   948 => x"486c87cc",
   949 => x"a6c49873",
   950 => x"05987058",
   951 => x"7cc487f4",
   952 => x"c348d4ff",
   953 => x"486c78ff",
   954 => x"a6c49873",
   955 => x"02987058",
   956 => x"486c87cc",
   957 => x"a6c49873",
   958 => x"05987058",
   959 => x"7cc587f4",
   960 => x"c148d4ff",
   961 => x"78c178d3",
   962 => x"9873486c",
   963 => x"7058a6c4",
   964 => x"87cc0298",
   965 => x"9873486c",
   966 => x"7058a6c4",
   967 => x"87f40598",
   968 => x"9d757cc4",
   969 => x"87d0c202",
   970 => x"7ed0d8c2",
   971 => x"ece5c21e",
   972 => x"87f8ea49",
   973 => x"987086c4",
   974 => x"c087c505",
   975 => x"87fcc248",
   976 => x"adb7c0c8",
   977 => x"4a87c404",
   978 => x"7587c48d",
   979 => x"6c4dc04a",
   980 => x"c8987348",
   981 => x"987058a6",
   982 => x"6c87cc02",
   983 => x"c8987348",
   984 => x"987058a6",
   985 => x"cd87f405",
   986 => x"48d4ff7c",
   987 => x"7278d4c1",
   988 => x"718ac149",
   989 => x"87d90299",
   990 => x"48bf976e",
   991 => x"7808d4ff",
   992 => x"80c1486e",
   993 => x"7258a6c4",
   994 => x"718ac149",
   995 => x"e7ff0599",
   996 => x"73486c87",
   997 => x"58a6c498",
   998 => x"cc029870",
   999 => x"73486c87",
  1000 => x"58a6c498",
  1001 => x"f4059870",
  1002 => x"c27cc487",
  1003 => x"e849ece5",
  1004 => x"9d7587d7",
  1005 => x"87f0fd05",
  1006 => x"9873486c",
  1007 => x"7058a6c4",
  1008 => x"87cd0298",
  1009 => x"9873486c",
  1010 => x"7058a6c4",
  1011 => x"f3ff0598",
  1012 => x"ff7cc587",
  1013 => x"d3c148d4",
  1014 => x"6c78c078",
  1015 => x"c4987348",
  1016 => x"987058a6",
  1017 => x"6c87cd02",
  1018 => x"c4987348",
  1019 => x"987058a6",
  1020 => x"87f3ff05",
  1021 => x"48c17cc4",
  1022 => x"48c087c2",
  1023 => x"cbf48ef4",
  1024 => x"5b5e0e87",
  1025 => x"1e0e5d5c",
  1026 => x"4cc04b71",
  1027 => x"04abb74d",
  1028 => x"c087e9c0",
  1029 => x"751ec3f5",
  1030 => x"87c4029d",
  1031 => x"87c24ac0",
  1032 => x"49724ac1",
  1033 => x"c487c2ea",
  1034 => x"c158a686",
  1035 => x"c2056e84",
  1036 => x"c14c7387",
  1037 => x"acb77385",
  1038 => x"87d7ff06",
  1039 => x"f326486e",
  1040 => x"5e0e87ca",
  1041 => x"0e5d5c5b",
  1042 => x"494c711e",
  1043 => x"bffce5c2",
  1044 => x"87edfe81",
  1045 => x"029d4d70",
  1046 => x"c287fcc0",
  1047 => x"754be0e0",
  1048 => x"ff49cb4a",
  1049 => x"7487c9c1",
  1050 => x"c291de49",
  1051 => x"7148d0e6",
  1052 => x"58a6c480",
  1053 => x"48e7c2c1",
  1054 => x"a1c8496e",
  1055 => x"7141204a",
  1056 => x"87f905aa",
  1057 => x"51105110",
  1058 => x"49745110",
  1059 => x"87eec5c1",
  1060 => x"49e0e0c2",
  1061 => x"c187c9f7",
  1062 => x"c149e0e4",
  1063 => x"c187f6c7",
  1064 => x"2687d2c8",
  1065 => x"4c87e5f1",
  1066 => x"6964616f",
  1067 => x"2e2e676e",
  1068 => x"2080002e",
  1069 => x"6b636142",
  1070 => x"616f4c00",
  1071 => x"2e2a2064",
  1072 => x"203a0020",
  1073 => x"42208000",
  1074 => x"006b6361",
  1075 => x"78452080",
  1076 => x"53007469",
  1077 => x"6e492044",
  1078 => x"2e2e7469",
  1079 => x"004b4f00",
  1080 => x"544f4f42",
  1081 => x"20202020",
  1082 => x"004d4f52",
  1083 => x"711e731e",
  1084 => x"e5c2494b",
  1085 => x"fc81bffc",
  1086 => x"4a7087c7",
  1087 => x"87c4029a",
  1088 => x"87e2e449",
  1089 => x"48fce5c2",
  1090 => x"497378c0",
  1091 => x"ef87e9c1",
  1092 => x"731e87fe",
  1093 => x"c44b711e",
  1094 => x"c1024aa3",
  1095 => x"8ac187c8",
  1096 => x"8a87dc02",
  1097 => x"87f1c002",
  1098 => x"c4c1058a",
  1099 => x"fce5c287",
  1100 => x"fcc002bf",
  1101 => x"88c14887",
  1102 => x"58c0e6c2",
  1103 => x"c287f2c0",
  1104 => x"49bffce5",
  1105 => x"e6c289d0",
  1106 => x"b7c059c0",
  1107 => x"e0c003a9",
  1108 => x"fce5c287",
  1109 => x"d878c048",
  1110 => x"fce5c287",
  1111 => x"80c148bf",
  1112 => x"58c0e6c2",
  1113 => x"e5c287cb",
  1114 => x"d048bffc",
  1115 => x"c0e6c280",
  1116 => x"c3497358",
  1117 => x"87d8ee87",
  1118 => x"5c5b5e0e",
  1119 => x"86f00e5d",
  1120 => x"c259a6d0",
  1121 => x"c04dd0d8",
  1122 => x"48a6c44c",
  1123 => x"e5c278c0",
  1124 => x"c048bffc",
  1125 => x"c106a8b7",
  1126 => x"d8c287c1",
  1127 => x"029848d0",
  1128 => x"c087f8c0",
  1129 => x"c81ec3f5",
  1130 => x"87c70266",
  1131 => x"c048a6c4",
  1132 => x"c487c578",
  1133 => x"78c148a6",
  1134 => x"e34966c4",
  1135 => x"86c487eb",
  1136 => x"84c14d70",
  1137 => x"c14866c4",
  1138 => x"58a6c880",
  1139 => x"bffce5c2",
  1140 => x"c603acb7",
  1141 => x"059d7587",
  1142 => x"c087c8ff",
  1143 => x"029d754c",
  1144 => x"c087e3c3",
  1145 => x"c81ec3f5",
  1146 => x"87c70266",
  1147 => x"c048a6cc",
  1148 => x"cc87c578",
  1149 => x"78c148a6",
  1150 => x"e24966cc",
  1151 => x"86c487eb",
  1152 => x"026e58a6",
  1153 => x"4987ebc2",
  1154 => x"699781cb",
  1155 => x"0299d049",
  1156 => x"c187d9c1",
  1157 => x"744becc3",
  1158 => x"c191cc49",
  1159 => x"c881e0e4",
  1160 => x"7a734aa1",
  1161 => x"ffc381c1",
  1162 => x"de497451",
  1163 => x"d0e6c291",
  1164 => x"c285714d",
  1165 => x"c17d97c1",
  1166 => x"e0c049a5",
  1167 => x"e0e0c251",
  1168 => x"d202bf97",
  1169 => x"c284c187",
  1170 => x"e0c24ba5",
  1171 => x"49db4ae0",
  1172 => x"87dcf9fe",
  1173 => x"cd87dbc1",
  1174 => x"51c049a5",
  1175 => x"a5c284c1",
  1176 => x"cb4a6e4b",
  1177 => x"c7f9fe49",
  1178 => x"87c6c187",
  1179 => x"91cc4974",
  1180 => x"81e0e4c1",
  1181 => x"c1c181c8",
  1182 => x"e0c279c2",
  1183 => x"02bf97e0",
  1184 => x"497487d8",
  1185 => x"84c191de",
  1186 => x"4bd0e6c2",
  1187 => x"e0c28371",
  1188 => x"49dd4ae0",
  1189 => x"87d8f8fe",
  1190 => x"4b7487d8",
  1191 => x"e6c293de",
  1192 => x"a3cb83d0",
  1193 => x"c151c049",
  1194 => x"4a6e7384",
  1195 => x"f7fe49cb",
  1196 => x"66c487fe",
  1197 => x"c880c148",
  1198 => x"b7c758a6",
  1199 => x"c5c003ac",
  1200 => x"fc056e87",
  1201 => x"b7c787dd",
  1202 => x"d3c003ac",
  1203 => x"de497487",
  1204 => x"d0e6c291",
  1205 => x"c151c081",
  1206 => x"acb7c784",
  1207 => x"87edff04",
  1208 => x"48f5e5c1",
  1209 => x"e5c150c0",
  1210 => x"50c248f4",
  1211 => x"48fce5c1",
  1212 => x"78deccc1",
  1213 => x"48f8e5c1",
  1214 => x"78f2c2c1",
  1215 => x"48c8e6c1",
  1216 => x"78d2c4c1",
  1217 => x"c04966cc",
  1218 => x"f087f3fb",
  1219 => x"87fce78e",
  1220 => x"c24a711e",
  1221 => x"725aece5",
  1222 => x"87dcf949",
  1223 => x"711e4f26",
  1224 => x"91cc494a",
  1225 => x"81e0e4c1",
  1226 => x"481181c1",
  1227 => x"58e8e5c2",
  1228 => x"49a2f0c0",
  1229 => x"87c8f6fe",
  1230 => x"ddd549c0",
  1231 => x"0e4f2687",
  1232 => x"5d5c5b5e",
  1233 => x"7186f00e",
  1234 => x"91cc494c",
  1235 => x"81e0e4c1",
  1236 => x"c47ea1c3",
  1237 => x"e5c248a6",
  1238 => x"6e78bfe0",
  1239 => x"c44abf97",
  1240 => x"2b724b66",
  1241 => x"124aa1c1",
  1242 => x"58a6cc48",
  1243 => x"83c19b70",
  1244 => x"699781c2",
  1245 => x"04abb749",
  1246 => x"4bc087c2",
  1247 => x"4abf976e",
  1248 => x"724966c8",
  1249 => x"c4b9ff31",
  1250 => x"4d739966",
  1251 => x"b5713572",
  1252 => x"5de4e5c2",
  1253 => x"c348d4ff",
  1254 => x"d0ff78ff",
  1255 => x"c0c848bf",
  1256 => x"a6d098c0",
  1257 => x"02987058",
  1258 => x"d0ff87d0",
  1259 => x"c0c848bf",
  1260 => x"a6c498c0",
  1261 => x"05987058",
  1262 => x"d0ff87f0",
  1263 => x"78e1c048",
  1264 => x"de48d4ff",
  1265 => x"7d0d7078",
  1266 => x"c848750d",
  1267 => x"d4ff28b7",
  1268 => x"48757808",
  1269 => x"ff28b7d0",
  1270 => x"757808d4",
  1271 => x"28b7d848",
  1272 => x"7808d4ff",
  1273 => x"48bfd0ff",
  1274 => x"98c0c0c8",
  1275 => x"7058a6c4",
  1276 => x"87d00298",
  1277 => x"48bfd0ff",
  1278 => x"98c0c0c8",
  1279 => x"7058a6c4",
  1280 => x"87f00598",
  1281 => x"c048d0ff",
  1282 => x"1ec778e0",
  1283 => x"e4c11ec0",
  1284 => x"e5c21ee0",
  1285 => x"c149bfe4",
  1286 => x"497487e1",
  1287 => x"87def7c0",
  1288 => x"e7e38ee4",
  1289 => x"1e731e87",
  1290 => x"fc494b71",
  1291 => x"497387d1",
  1292 => x"e387ccfc",
  1293 => x"731e87da",
  1294 => x"c24b711e",
  1295 => x"d5024aa3",
  1296 => x"058ac187",
  1297 => x"e5c287db",
  1298 => x"d402bff8",
  1299 => x"88c14887",
  1300 => x"58fce5c2",
  1301 => x"e5c287cb",
  1302 => x"c148bff8",
  1303 => x"fce5c280",
  1304 => x"c01ec758",
  1305 => x"e0e4c11e",
  1306 => x"e4e5c21e",
  1307 => x"87cb49bf",
  1308 => x"f6c04973",
  1309 => x"8ef487c8",
  1310 => x"0e87d5e2",
  1311 => x"5d5c5b5e",
  1312 => x"86d8ff0e",
  1313 => x"c859a6dc",
  1314 => x"78c048a6",
  1315 => x"78c080c4",
  1316 => x"c280c44d",
  1317 => x"78bff8e5",
  1318 => x"c348d4ff",
  1319 => x"d0ff78ff",
  1320 => x"c0c848bf",
  1321 => x"a6c498c0",
  1322 => x"02987058",
  1323 => x"d0ff87d0",
  1324 => x"c0c848bf",
  1325 => x"a6c498c0",
  1326 => x"05987058",
  1327 => x"d0ff87f0",
  1328 => x"78e1c048",
  1329 => x"d448d4ff",
  1330 => x"f6deff78",
  1331 => x"48d4ff87",
  1332 => x"d478ffc3",
  1333 => x"d4ff48a6",
  1334 => x"66d478bf",
  1335 => x"a8fbc048",
  1336 => x"87d3c102",
  1337 => x"4a66f8c0",
  1338 => x"7e6a82c4",
  1339 => x"c2c11e72",
  1340 => x"66c448f9",
  1341 => x"4aa1c849",
  1342 => x"aa714120",
  1343 => x"1087f905",
  1344 => x"c04a2651",
  1345 => x"c84966f8",
  1346 => x"d0ccc181",
  1347 => x"c7496a79",
  1348 => x"5166d481",
  1349 => x"1ed81ec1",
  1350 => x"81c8496a",
  1351 => x"87faddff",
  1352 => x"66d086c8",
  1353 => x"a8b7c048",
  1354 => x"c187c401",
  1355 => x"d087c84d",
  1356 => x"88c14866",
  1357 => x"d458a6d4",
  1358 => x"f4ca0266",
  1359 => x"66c0c187",
  1360 => x"ca03adb7",
  1361 => x"d4ff87eb",
  1362 => x"78ffc348",
  1363 => x"ff48a6d4",
  1364 => x"d478bfd4",
  1365 => x"c6c14866",
  1366 => x"58a6c488",
  1367 => x"c0029870",
  1368 => x"c94887e6",
  1369 => x"58a6c488",
  1370 => x"c4029870",
  1371 => x"c14887d5",
  1372 => x"58a6c488",
  1373 => x"c1029870",
  1374 => x"c44887e3",
  1375 => x"7058a688",
  1376 => x"fec30298",
  1377 => x"87d3c987",
  1378 => x"c10566d8",
  1379 => x"d4ff87c5",
  1380 => x"78ffc348",
  1381 => x"1eca1ec0",
  1382 => x"93cc4b75",
  1383 => x"8366c0c1",
  1384 => x"6c4ca3c4",
  1385 => x"f1dbff49",
  1386 => x"de1ec187",
  1387 => x"ff496c1e",
  1388 => x"d087e7db",
  1389 => x"49a3c886",
  1390 => x"79d0ccc1",
  1391 => x"adb766d0",
  1392 => x"c187c504",
  1393 => x"87dac885",
  1394 => x"c14866d0",
  1395 => x"58a6d488",
  1396 => x"ff87cfc8",
  1397 => x"d887ecda",
  1398 => x"c5c858a6",
  1399 => x"f3dcff87",
  1400 => x"58a6cc87",
  1401 => x"a8b766cc",
  1402 => x"cc87c606",
  1403 => x"66c848a6",
  1404 => x"dfdcff78",
  1405 => x"a8ecc087",
  1406 => x"87c7c205",
  1407 => x"c10566d8",
  1408 => x"497587f7",
  1409 => x"f8c091cc",
  1410 => x"a1c48166",
  1411 => x"c14c6a4a",
  1412 => x"66c84aa1",
  1413 => x"7997c252",
  1414 => x"ccc181c8",
  1415 => x"d4ff79de",
  1416 => x"78ffc348",
  1417 => x"ff48a6d4",
  1418 => x"d478bfd4",
  1419 => x"e8c00266",
  1420 => x"fbc04887",
  1421 => x"e0c002a8",
  1422 => x"9766d487",
  1423 => x"ff84c17c",
  1424 => x"ffc348d4",
  1425 => x"48a6d478",
  1426 => x"78bfd4ff",
  1427 => x"c80266d4",
  1428 => x"fbc04887",
  1429 => x"e0ff05a8",
  1430 => x"54e0c087",
  1431 => x"c054c1c2",
  1432 => x"66d07c97",
  1433 => x"c504adb7",
  1434 => x"c585c187",
  1435 => x"66d087f4",
  1436 => x"d488c148",
  1437 => x"e9c558a6",
  1438 => x"c6d8ff87",
  1439 => x"58a6d887",
  1440 => x"c887dfc5",
  1441 => x"66d84866",
  1442 => x"c4c505a8",
  1443 => x"48a6dc87",
  1444 => x"d9ff78c0",
  1445 => x"a6d887fe",
  1446 => x"f7d9ff58",
  1447 => x"a6e4c087",
  1448 => x"a8ecc058",
  1449 => x"87cac005",
  1450 => x"48a6e0c0",
  1451 => x"c07866d4",
  1452 => x"d4ff87c6",
  1453 => x"78ffc348",
  1454 => x"91cc4975",
  1455 => x"4866f8c0",
  1456 => x"a6c48071",
  1457 => x"c3496e58",
  1458 => x"5166d481",
  1459 => x"4966e0c0",
  1460 => x"66d481c1",
  1461 => x"7148c189",
  1462 => x"c1497030",
  1463 => x"c14a6e89",
  1464 => x"97097282",
  1465 => x"486e0979",
  1466 => x"e5c250c2",
  1467 => x"d449bfe0",
  1468 => x"9729b766",
  1469 => x"71484a6a",
  1470 => x"a6e8c098",
  1471 => x"c4486e58",
  1472 => x"58a6c880",
  1473 => x"4cbf66c4",
  1474 => x"c84866d8",
  1475 => x"c002a866",
  1476 => x"e0c087c9",
  1477 => x"78c048a6",
  1478 => x"c087c6c0",
  1479 => x"c148a6e0",
  1480 => x"66e0c078",
  1481 => x"1ee0c01e",
  1482 => x"d5ff4974",
  1483 => x"86c887ec",
  1484 => x"c058a6d8",
  1485 => x"c106a8b7",
  1486 => x"66d487da",
  1487 => x"bf66c484",
  1488 => x"81e0c049",
  1489 => x"c14b8974",
  1490 => x"714ac2c3",
  1491 => x"87e0e5fe",
  1492 => x"66dc84c2",
  1493 => x"c080c148",
  1494 => x"c058a6e0",
  1495 => x"c14966e4",
  1496 => x"02a97081",
  1497 => x"c087c9c0",
  1498 => x"c048a6e0",
  1499 => x"87c6c078",
  1500 => x"48a6e0c0",
  1501 => x"e0c078c1",
  1502 => x"66c81e66",
  1503 => x"e0c049bf",
  1504 => x"71897481",
  1505 => x"ff49741e",
  1506 => x"c887cfd4",
  1507 => x"a8b7c086",
  1508 => x"87fefe01",
  1509 => x"c00266dc",
  1510 => x"496e87d2",
  1511 => x"66dc81c2",
  1512 => x"c8496e51",
  1513 => x"ffccc181",
  1514 => x"87cdc079",
  1515 => x"81c2496e",
  1516 => x"c8496e51",
  1517 => x"e5d0c181",
  1518 => x"b766d079",
  1519 => x"c5c004ad",
  1520 => x"c085c187",
  1521 => x"66d087dc",
  1522 => x"d488c148",
  1523 => x"d1c058a6",
  1524 => x"eed2ff87",
  1525 => x"58a6d887",
  1526 => x"ff87c7c0",
  1527 => x"d887e4d2",
  1528 => x"66d458a6",
  1529 => x"87c9c002",
  1530 => x"b766c0c1",
  1531 => x"d5f504ad",
  1532 => x"adb7c787",
  1533 => x"87dcc003",
  1534 => x"91cc4975",
  1535 => x"8166f8c0",
  1536 => x"6a4aa1c4",
  1537 => x"c852c04a",
  1538 => x"c179c081",
  1539 => x"adb7c785",
  1540 => x"87e4ff04",
  1541 => x"c00266d8",
  1542 => x"f8c087eb",
  1543 => x"d4c14966",
  1544 => x"66f8c081",
  1545 => x"82d5c14a",
  1546 => x"51c252c0",
  1547 => x"4966f8c0",
  1548 => x"c181dcc1",
  1549 => x"c079decc",
  1550 => x"c14966f8",
  1551 => x"c3c181d8",
  1552 => x"d6c079c5",
  1553 => x"66f8c087",
  1554 => x"81d8c149",
  1555 => x"79ccc3c1",
  1556 => x"4966f8c0",
  1557 => x"c281dcc1",
  1558 => x"c179f5ca",
  1559 => x"c04af6d0",
  1560 => x"c14966f8",
  1561 => x"797281e8",
  1562 => x"48bfd0ff",
  1563 => x"98c0c0c8",
  1564 => x"7058a6c4",
  1565 => x"d1c00298",
  1566 => x"bfd0ff87",
  1567 => x"c0c0c848",
  1568 => x"58a6c498",
  1569 => x"ff059870",
  1570 => x"d0ff87ef",
  1571 => x"78e0c048",
  1572 => x"ff4866cc",
  1573 => x"d1ff8ed8",
  1574 => x"c71e87f2",
  1575 => x"c11ec01e",
  1576 => x"c21ee0e4",
  1577 => x"49bfe4e5",
  1578 => x"c187d0ef",
  1579 => x"c049e0e4",
  1580 => x"f487e2e7",
  1581 => x"1e4f268e",
  1582 => x"c287c6ca",
  1583 => x"c048c0e6",
  1584 => x"48d4ff50",
  1585 => x"c178ffc3",
  1586 => x"fe49d3c3",
  1587 => x"fe87fdde",
  1588 => x"7087c8e8",
  1589 => x"87cd0298",
  1590 => x"87c5f4fe",
  1591 => x"c4029870",
  1592 => x"c24ac187",
  1593 => x"724ac087",
  1594 => x"87c8029a",
  1595 => x"49ddc3c1",
  1596 => x"87d8defe",
  1597 => x"bfd0d7c2",
  1598 => x"e3d5ff49",
  1599 => x"f8e5c287",
  1600 => x"c278c048",
  1601 => x"c048e4e5",
  1602 => x"cdfe4978",
  1603 => x"87ddc387",
  1604 => x"c087c2c9",
  1605 => x"ff87ede6",
  1606 => x"4f2687f6",
  1607 => x"000010e0",
  1608 => x"00000002",
  1609 => x"00002990",
  1610 => x"00001042",
  1611 => x"00000002",
  1612 => x"000029ae",
  1613 => x"00001042",
  1614 => x"00000002",
  1615 => x"000029cc",
  1616 => x"00001042",
  1617 => x"00000002",
  1618 => x"000029ea",
  1619 => x"00001042",
  1620 => x"00000002",
  1621 => x"00002a08",
  1622 => x"00001042",
  1623 => x"00000002",
  1624 => x"00002a26",
  1625 => x"00001042",
  1626 => x"00000002",
  1627 => x"00002a44",
  1628 => x"00001042",
  1629 => x"00000002",
  1630 => x"00000000",
  1631 => x"0000131e",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"00001112",
  1635 => x"d5c11e1e",
  1636 => x"58a6c487",
  1637 => x"1e4f2626",
  1638 => x"f0fe4a71",
  1639 => x"cd78c048",
  1640 => x"c10a7a0a",
  1641 => x"fe49ede6",
  1642 => x"2687e1db",
  1643 => x"7465534f",
  1644 => x"6e616820",
  1645 => x"72656c64",
  1646 => x"6e49000a",
  1647 => x"746e6920",
  1648 => x"75727265",
  1649 => x"63207470",
  1650 => x"74736e6f",
  1651 => x"74637572",
  1652 => x"000a726f",
  1653 => x"fae6c11e",
  1654 => x"efdafe49",
  1655 => x"cce6c187",
  1656 => x"87f3fe49",
  1657 => x"fe1e4f26",
  1658 => x"2648bff0",
  1659 => x"f0fe1e4f",
  1660 => x"2678c148",
  1661 => x"f0fe1e4f",
  1662 => x"2678c048",
  1663 => x"4a711e4f",
  1664 => x"a2c47ac0",
  1665 => x"c879c049",
  1666 => x"79c049a2",
  1667 => x"c049a2cc",
  1668 => x"0e4f2679",
  1669 => x"0e5c5b5e",
  1670 => x"4c7186f8",
  1671 => x"cc49a4c8",
  1672 => x"486b4ba4",
  1673 => x"a6c480c1",
  1674 => x"c898cf58",
  1675 => x"486958a6",
  1676 => x"05a866c4",
  1677 => x"486b87d4",
  1678 => x"a6c480c1",
  1679 => x"c898cf58",
  1680 => x"486958a6",
  1681 => x"02a866c4",
  1682 => x"e8fe87ec",
  1683 => x"a4d0c187",
  1684 => x"c4486b49",
  1685 => x"58a6c490",
  1686 => x"66d48170",
  1687 => x"c1486b79",
  1688 => x"58a6c880",
  1689 => x"7b7098cf",
  1690 => x"fd87d2c1",
  1691 => x"8ef887ff",
  1692 => x"4d2687c2",
  1693 => x"4b264c26",
  1694 => x"5e0e4f26",
  1695 => x"0e5d5c5b",
  1696 => x"4d7186f8",
  1697 => x"6d4ca5c4",
  1698 => x"05a86c48",
  1699 => x"48ff87c5",
  1700 => x"fd87e5c0",
  1701 => x"a5d087df",
  1702 => x"c4486c4b",
  1703 => x"58a6c490",
  1704 => x"4b6b8370",
  1705 => x"6c9bffc3",
  1706 => x"c880c148",
  1707 => x"98cf58a6",
  1708 => x"f8fc7c70",
  1709 => x"48497387",
  1710 => x"f5fe8ef8",
  1711 => x"1e731e87",
  1712 => x"f0fc86f8",
  1713 => x"4bbfe087",
  1714 => x"c0e0c049",
  1715 => x"e7c00299",
  1716 => x"c34a7387",
  1717 => x"e9c29aff",
  1718 => x"c448bfe2",
  1719 => x"58a6c490",
  1720 => x"49f2e9c2",
  1721 => x"79728170",
  1722 => x"bfe2e9c2",
  1723 => x"c880c148",
  1724 => x"98cf58a6",
  1725 => x"58e6e9c2",
  1726 => x"c0d04973",
  1727 => x"f2c00299",
  1728 => x"eae9c287",
  1729 => x"e9c248bf",
  1730 => x"02a8bfee",
  1731 => x"c287e4c0",
  1732 => x"48bfeae9",
  1733 => x"a6c490c4",
  1734 => x"f2eac258",
  1735 => x"e0817049",
  1736 => x"c2786948",
  1737 => x"48bfeae9",
  1738 => x"a6c880c1",
  1739 => x"c298cf58",
  1740 => x"fa58eee9",
  1741 => x"a6c487f0",
  1742 => x"87f1fa58",
  1743 => x"f5fc8ef8",
  1744 => x"e9c21e87",
  1745 => x"f4fa49e2",
  1746 => x"fdeac187",
  1747 => x"87c7f949",
  1748 => x"2687f5c3",
  1749 => x"1e731e4f",
  1750 => x"49e2e9c2",
  1751 => x"7087dbfc",
  1752 => x"aab7c04a",
  1753 => x"87ccc204",
  1754 => x"05aaf0c3",
  1755 => x"f0c187c9",
  1756 => x"78c148c0",
  1757 => x"c387edc1",
  1758 => x"c905aae0",
  1759 => x"c4f0c187",
  1760 => x"c178c148",
  1761 => x"f0c187de",
  1762 => x"c602bfc4",
  1763 => x"a2c0c287",
  1764 => x"7287c24b",
  1765 => x"c0f0c14b",
  1766 => x"e0c002bf",
  1767 => x"c4497387",
  1768 => x"c19129b7",
  1769 => x"7381c8f0",
  1770 => x"c29acf4a",
  1771 => x"7248c192",
  1772 => x"ff4a7030",
  1773 => x"694872ba",
  1774 => x"db797098",
  1775 => x"c4497387",
  1776 => x"c19129b7",
  1777 => x"7381c8f0",
  1778 => x"c29acf4a",
  1779 => x"7248c392",
  1780 => x"484a7030",
  1781 => x"7970b069",
  1782 => x"48c4f0c1",
  1783 => x"f0c178c0",
  1784 => x"78c048c0",
  1785 => x"49e2e9c2",
  1786 => x"7087cffa",
  1787 => x"aab7c04a",
  1788 => x"87f4fd03",
  1789 => x"87c448c0",
  1790 => x"4c264d26",
  1791 => x"4f264b26",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000000",
  1807 => x"00000000",
  1808 => x"00000000",
  1809 => x"00000000",
  1810 => x"724ac01e",
  1811 => x"c191c449",
  1812 => x"c081c8f0",
  1813 => x"d082c179",
  1814 => x"ee04aab7",
  1815 => x"0e4f2687",
  1816 => x"5d5c5b5e",
  1817 => x"f64d710e",
  1818 => x"4a7587cb",
  1819 => x"922ab7c4",
  1820 => x"82c8f0c1",
  1821 => x"9ccf4c75",
  1822 => x"496a94c2",
  1823 => x"c32b744b",
  1824 => x"7448c29b",
  1825 => x"ff4c7030",
  1826 => x"714874bc",
  1827 => x"f57a7098",
  1828 => x"487387db",
  1829 => x"1e87e1fd",
  1830 => x"bfd0ff1e",
  1831 => x"c0c0c848",
  1832 => x"58a6c498",
  1833 => x"d0029870",
  1834 => x"bfd0ff87",
  1835 => x"c0c0c848",
  1836 => x"58a6c498",
  1837 => x"f0059870",
  1838 => x"48d0ff87",
  1839 => x"7178e1c4",
  1840 => x"08d4ff48",
  1841 => x"4866c878",
  1842 => x"7808d4ff",
  1843 => x"1e4f2626",
  1844 => x"c84a711e",
  1845 => x"721e4966",
  1846 => x"87fbfe49",
  1847 => x"d0ff86c4",
  1848 => x"c0c848bf",
  1849 => x"a6c498c0",
  1850 => x"02987058",
  1851 => x"d0ff87d0",
  1852 => x"c0c848bf",
  1853 => x"a6c498c0",
  1854 => x"05987058",
  1855 => x"d0ff87f0",
  1856 => x"78e0c048",
  1857 => x"1e4f2626",
  1858 => x"4b711e73",
  1859 => x"731e66c8",
  1860 => x"a2e0c14a",
  1861 => x"87f7fe49",
  1862 => x"2687c426",
  1863 => x"264c264d",
  1864 => x"1e4f264b",
  1865 => x"bfd0ff1e",
  1866 => x"c0c0c848",
  1867 => x"58a6c498",
  1868 => x"d0029870",
  1869 => x"bfd0ff87",
  1870 => x"c0c0c848",
  1871 => x"58a6c498",
  1872 => x"f0059870",
  1873 => x"48d0ff87",
  1874 => x"7178c9c4",
  1875 => x"08d4ff48",
  1876 => x"4f262678",
  1877 => x"4a711e1e",
  1878 => x"87c7ff49",
  1879 => x"48bfd0ff",
  1880 => x"98c0c0c8",
  1881 => x"7058a6c4",
  1882 => x"87d00298",
  1883 => x"48bfd0ff",
  1884 => x"98c0c0c8",
  1885 => x"7058a6c4",
  1886 => x"87f00598",
  1887 => x"c848d0ff",
  1888 => x"4f262678",
  1889 => x"1e1e731e",
  1890 => x"ebc24b71",
  1891 => x"c302bffe",
  1892 => x"87ccc387",
  1893 => x"48bfd0ff",
  1894 => x"98c0c0c8",
  1895 => x"7058a6c4",
  1896 => x"87d00298",
  1897 => x"48bfd0ff",
  1898 => x"98c0c0c8",
  1899 => x"7058a6c4",
  1900 => x"87f00598",
  1901 => x"c448d0ff",
  1902 => x"487378c9",
  1903 => x"ffb0e0c0",
  1904 => x"c27808d4",
  1905 => x"c048f2eb",
  1906 => x"0266cc78",
  1907 => x"ffc387c5",
  1908 => x"c087c249",
  1909 => x"faebc249",
  1910 => x"0266d059",
  1911 => x"d5c587c6",
  1912 => x"87c44ad5",
  1913 => x"4affffcf",
  1914 => x"5afeebc2",
  1915 => x"48feebc2",
  1916 => x"c42678c1",
  1917 => x"264d2687",
  1918 => x"264b264c",
  1919 => x"5b5e0e4f",
  1920 => x"710e5d5c",
  1921 => x"faebc24a",
  1922 => x"9a724cbf",
  1923 => x"4987cb02",
  1924 => x"f6c191c8",
  1925 => x"83714bfe",
  1926 => x"fac187c4",
  1927 => x"4dc04bfe",
  1928 => x"99744913",
  1929 => x"bff6ebc2",
  1930 => x"ffb87148",
  1931 => x"c17808d4",
  1932 => x"c8852cb7",
  1933 => x"e704adb7",
  1934 => x"f2ebc287",
  1935 => x"80c848bf",
  1936 => x"58f6ebc2",
  1937 => x"1e87eefe",
  1938 => x"4b711e73",
  1939 => x"029a4a13",
  1940 => x"497287cb",
  1941 => x"1387e6fe",
  1942 => x"f5059a4a",
  1943 => x"87d9fe87",
  1944 => x"ebc21e1e",
  1945 => x"c249bff2",
  1946 => x"c148f2eb",
  1947 => x"c0c478a1",
  1948 => x"db03a9b7",
  1949 => x"48d4ff87",
  1950 => x"bff6ebc2",
  1951 => x"f2ebc278",
  1952 => x"ebc249bf",
  1953 => x"a1c148f2",
  1954 => x"b7c0c478",
  1955 => x"87e504a9",
  1956 => x"48bfd0ff",
  1957 => x"98c0c0c8",
  1958 => x"7058a6c4",
  1959 => x"87d00298",
  1960 => x"48bfd0ff",
  1961 => x"98c0c0c8",
  1962 => x"7058a6c4",
  1963 => x"87f00598",
  1964 => x"c848d0ff",
  1965 => x"feebc278",
  1966 => x"2678c048",
  1967 => x"00004f26",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"005f5f00",
  1971 => x"03000000",
  1972 => x"03030003",
  1973 => x"7f140000",
  1974 => x"7f7f147f",
  1975 => x"24000014",
  1976 => x"3a6b6b2e",
  1977 => x"6a4c0012",
  1978 => x"566c1836",
  1979 => x"7e300032",
  1980 => x"3a77594f",
  1981 => x"00004068",
  1982 => x"00030704",
  1983 => x"00000000",
  1984 => x"41633e1c",
  1985 => x"00000000",
  1986 => x"1c3e6341",
  1987 => x"2a080000",
  1988 => x"3e1c1c3e",
  1989 => x"0800082a",
  1990 => x"083e3e08",
  1991 => x"00000008",
  1992 => x"0060e080",
  1993 => x"08000000",
  1994 => x"08080808",
  1995 => x"00000008",
  1996 => x"00606000",
  1997 => x"60400000",
  1998 => x"060c1830",
  1999 => x"3e000103",
  2000 => x"7f4d597f",
  2001 => x"0400003e",
  2002 => x"007f7f06",
  2003 => x"42000000",
  2004 => x"4f597163",
  2005 => x"22000046",
  2006 => x"7f494963",
  2007 => x"1c180036",
  2008 => x"7f7f1316",
  2009 => x"27000010",
  2010 => x"7d454567",
  2011 => x"3c000039",
  2012 => x"79494b7e",
  2013 => x"01000030",
  2014 => x"0f797101",
  2015 => x"36000007",
  2016 => x"7f49497f",
  2017 => x"06000036",
  2018 => x"3f69494f",
  2019 => x"0000001e",
  2020 => x"00666600",
  2021 => x"00000000",
  2022 => x"0066e680",
  2023 => x"08000000",
  2024 => x"22141408",
  2025 => x"14000022",
  2026 => x"14141414",
  2027 => x"22000014",
  2028 => x"08141422",
  2029 => x"02000008",
  2030 => x"0f595103",
  2031 => x"7f3e0006",
  2032 => x"1f555d41",
  2033 => x"7e00001e",
  2034 => x"7f09097f",
  2035 => x"7f00007e",
  2036 => x"7f49497f",
  2037 => x"1c000036",
  2038 => x"4141633e",
  2039 => x"7f000041",
  2040 => x"3e63417f",
  2041 => x"7f00001c",
  2042 => x"4149497f",
  2043 => x"7f000041",
  2044 => x"0109097f",
  2045 => x"3e000001",
  2046 => x"7b49417f",
  2047 => x"7f00007a",
  2048 => x"7f08087f",
  2049 => x"0000007f",
  2050 => x"417f7f41",
  2051 => x"20000000",
  2052 => x"7f404060",
  2053 => x"7f7f003f",
  2054 => x"63361c08",
  2055 => x"7f000041",
  2056 => x"4040407f",
  2057 => x"7f7f0040",
  2058 => x"7f060c06",
  2059 => x"7f7f007f",
  2060 => x"7f180c06",
  2061 => x"3e00007f",
  2062 => x"7f41417f",
  2063 => x"7f00003e",
  2064 => x"0f09097f",
  2065 => x"7f3e0006",
  2066 => x"7e7f6141",
  2067 => x"7f000040",
  2068 => x"7f19097f",
  2069 => x"26000066",
  2070 => x"7b594d6f",
  2071 => x"01000032",
  2072 => x"017f7f01",
  2073 => x"3f000001",
  2074 => x"7f40407f",
  2075 => x"0f00003f",
  2076 => x"3f70703f",
  2077 => x"7f7f000f",
  2078 => x"7f301830",
  2079 => x"6341007f",
  2080 => x"361c1c36",
  2081 => x"03014163",
  2082 => x"067c7c06",
  2083 => x"71610103",
  2084 => x"43474d59",
  2085 => x"00000041",
  2086 => x"41417f7f",
  2087 => x"03010000",
  2088 => x"30180c06",
  2089 => x"00004060",
  2090 => x"7f7f4141",
  2091 => x"0c080000",
  2092 => x"0c060306",
  2093 => x"80800008",
  2094 => x"80808080",
  2095 => x"00000080",
  2096 => x"04070300",
  2097 => x"20000000",
  2098 => x"7c545474",
  2099 => x"7f000078",
  2100 => x"7c44447f",
  2101 => x"38000038",
  2102 => x"4444447c",
  2103 => x"38000000",
  2104 => x"7f44447c",
  2105 => x"3800007f",
  2106 => x"5c54547c",
  2107 => x"04000018",
  2108 => x"05057f7e",
  2109 => x"18000000",
  2110 => x"fca4a4bc",
  2111 => x"7f00007c",
  2112 => x"7c04047f",
  2113 => x"00000078",
  2114 => x"407d3d00",
  2115 => x"80000000",
  2116 => x"7dfd8080",
  2117 => x"7f000000",
  2118 => x"6c38107f",
  2119 => x"00000044",
  2120 => x"407f3f00",
  2121 => x"7c7c0000",
  2122 => x"7c0c180c",
  2123 => x"7c000078",
  2124 => x"7c04047c",
  2125 => x"38000078",
  2126 => x"7c44447c",
  2127 => x"fc000038",
  2128 => x"3c2424fc",
  2129 => x"18000018",
  2130 => x"fc24243c",
  2131 => x"7c0000fc",
  2132 => x"0c04047c",
  2133 => x"48000008",
  2134 => x"7454545c",
  2135 => x"04000020",
  2136 => x"44447f3f",
  2137 => x"3c000000",
  2138 => x"7c40407c",
  2139 => x"1c00007c",
  2140 => x"3c60603c",
  2141 => x"7c3c001c",
  2142 => x"7c603060",
  2143 => x"6c44003c",
  2144 => x"6c381038",
  2145 => x"1c000044",
  2146 => x"3c60e0bc",
  2147 => x"4400001c",
  2148 => x"4c5c7464",
  2149 => x"08000044",
  2150 => x"41773e08",
  2151 => x"00000041",
  2152 => x"007f7f00",
  2153 => x"41000000",
  2154 => x"083e7741",
  2155 => x"01020008",
  2156 => x"02020301",
  2157 => x"7f7f0001",
  2158 => x"7f7f7f7f",
  2159 => x"0808007f",
  2160 => x"3e3e1c1c",
  2161 => x"7f7f7f7f",
  2162 => x"1c1c3e3e",
  2163 => x"10000808",
  2164 => x"187c7c18",
  2165 => x"10000010",
  2166 => x"307c7c30",
  2167 => x"30100010",
  2168 => x"1e786060",
  2169 => x"66420006",
  2170 => x"663c183c",
  2171 => x"38780042",
  2172 => x"6cc6c26a",
  2173 => x"00600038",
  2174 => x"00006000",
  2175 => x"5e0e0060",
  2176 => x"0e5d5c5b",
  2177 => x"c24c711e",
  2178 => x"4bbfc6ec",
  2179 => x"48caecc2",
  2180 => x"062778c0",
  2181 => x"bf00002b",
  2182 => x"9949bf97",
  2183 => x"87c8c102",
  2184 => x"ecc21ec0",
  2185 => x"744dbfca",
  2186 => x"87c702ad",
  2187 => x"c048a6c4",
  2188 => x"c487c578",
  2189 => x"78c148a6",
  2190 => x"751e66c4",
  2191 => x"87c4ed49",
  2192 => x"e0c086c8",
  2193 => x"87f5ee49",
  2194 => x"6a4aa3c4",
  2195 => x"87f7ef49",
  2196 => x"c287cdf0",
  2197 => x"48bfcaec",
  2198 => x"ecc280c1",
  2199 => x"83cc58ce",
  2200 => x"99496b97",
  2201 => x"87f8fe05",
  2202 => x"bfcaecc2",
  2203 => x"adb7c84d",
  2204 => x"c087d903",
  2205 => x"ecc21e1e",
  2206 => x"ec49bfca",
  2207 => x"86c887c6",
  2208 => x"c187ddef",
  2209 => x"adb7c885",
  2210 => x"87e7ff04",
  2211 => x"264d2626",
  2212 => x"264b264c",
  2213 => x"4a711e4f",
  2214 => x"5acaecc2",
  2215 => x"bfceecc2",
  2216 => x"87dafd49",
  2217 => x"bfcaecc2",
  2218 => x"c289c149",
  2219 => x"7159d2ec",
  2220 => x"2687cbfd",
  2221 => x"c0c11e4f",
  2222 => x"87d8ea49",
  2223 => x"48fbd6c2",
  2224 => x"4f2678c0",
  2225 => x"5c5b5e0e",
  2226 => x"86f40e5d",
  2227 => x"c048a6c8",
  2228 => x"7ebfec78",
  2229 => x"ecc280fc",
  2230 => x"c278bfc6",
  2231 => x"4dbfd2ec",
  2232 => x"c74cbfe8",
  2233 => x"87f7e549",
  2234 => x"99c24970",
  2235 => x"c287cf05",
  2236 => x"49bff3d6",
  2237 => x"996eb9ff",
  2238 => x"c00299c1",
  2239 => x"49c787ee",
  2240 => x"7087dce5",
  2241 => x"87cd0298",
  2242 => x"c787cae1",
  2243 => x"87cfe549",
  2244 => x"f3059870",
  2245 => x"fbd6c287",
  2246 => x"bac14abf",
  2247 => x"5affd6c2",
  2248 => x"49a2c0c1",
  2249 => x"c887ede8",
  2250 => x"78c148a6",
  2251 => x"48f3d6c2",
  2252 => x"d6c2786e",
  2253 => x"c105bffb",
  2254 => x"a6c487da",
  2255 => x"c0c0c848",
  2256 => x"ffd6c278",
  2257 => x"bf976e7e",
  2258 => x"c1486e49",
  2259 => x"58a6c480",
  2260 => x"87cbe471",
  2261 => x"c3029870",
  2262 => x"b466c487",
  2263 => x"c14866c4",
  2264 => x"a6c828b7",
  2265 => x"05987058",
  2266 => x"7487daff",
  2267 => x"99ffc349",
  2268 => x"49c01e71",
  2269 => x"7487d0e6",
  2270 => x"29b7c849",
  2271 => x"49c11e71",
  2272 => x"c887c4e6",
  2273 => x"49fdc386",
  2274 => x"c387d4e3",
  2275 => x"cee349fa",
  2276 => x"87cac887",
  2277 => x"ffc34974",
  2278 => x"2cb7c899",
  2279 => x"9c74b471",
  2280 => x"ff87dd02",
  2281 => x"6e7ebfc8",
  2282 => x"f7d6c249",
  2283 => x"c0c289bf",
  2284 => x"87c403a9",
  2285 => x"87ce4cc0",
  2286 => x"48f7d6c2",
  2287 => x"87c6786e",
  2288 => x"48f7d6c2",
  2289 => x"497478c0",
  2290 => x"ce0599c8",
  2291 => x"49f5c387",
  2292 => x"7087cce2",
  2293 => x"0299c249",
  2294 => x"c287edc0",
  2295 => x"02bfceec",
  2296 => x"c14887c9",
  2297 => x"d2ecc288",
  2298 => x"c287d858",
  2299 => x"49bfcaec",
  2300 => x"66c491cc",
  2301 => x"7ea1c881",
  2302 => x"c002bf6e",
  2303 => x"ff4b87c5",
  2304 => x"c80f7349",
  2305 => x"78c148a6",
  2306 => x"99c44974",
  2307 => x"c387ce05",
  2308 => x"cae149f2",
  2309 => x"c2497087",
  2310 => x"fdc00299",
  2311 => x"48a6c887",
  2312 => x"bfcaecc2",
  2313 => x"4966c878",
  2314 => x"ecc289c1",
  2315 => x"6e7ebfce",
  2316 => x"c006a9b7",
  2317 => x"c14887c9",
  2318 => x"d2ecc280",
  2319 => x"c887d658",
  2320 => x"91cc4966",
  2321 => x"c88166c4",
  2322 => x"bf6e7ea1",
  2323 => x"87c5c002",
  2324 => x"7349fe4b",
  2325 => x"48a6c80f",
  2326 => x"fdc378c1",
  2327 => x"fedfff49",
  2328 => x"c2497087",
  2329 => x"eec00299",
  2330 => x"ceecc287",
  2331 => x"c9c002bf",
  2332 => x"ceecc287",
  2333 => x"c078c048",
  2334 => x"ecc287d8",
  2335 => x"cc49bfca",
  2336 => x"8166c491",
  2337 => x"6e7ea1c8",
  2338 => x"c5c002bf",
  2339 => x"49fd4b87",
  2340 => x"a6c80f73",
  2341 => x"c378c148",
  2342 => x"dfff49fa",
  2343 => x"497087c1",
  2344 => x"c10299c2",
  2345 => x"a6c887c0",
  2346 => x"caecc248",
  2347 => x"66c878bf",
  2348 => x"c488c148",
  2349 => x"ecc258a6",
  2350 => x"6e48bfce",
  2351 => x"c003a8b7",
  2352 => x"ecc287c9",
  2353 => x"786e48ce",
  2354 => x"c887d6c0",
  2355 => x"91cc4966",
  2356 => x"c88166c4",
  2357 => x"bf6e7ea1",
  2358 => x"87c5c002",
  2359 => x"7349fc4b",
  2360 => x"48a6c80f",
  2361 => x"ecc278c1",
  2362 => x"c04abfce",
  2363 => x"c006aab7",
  2364 => x"8ac187c9",
  2365 => x"01aab7c0",
  2366 => x"7487f7ff",
  2367 => x"99f0c349",
  2368 => x"87cfc005",
  2369 => x"ff49dac1",
  2370 => x"7087d4dd",
  2371 => x"0299c249",
  2372 => x"c287cec1",
  2373 => x"7ebfc6ec",
  2374 => x"c248a6c4",
  2375 => x"78bfceec",
  2376 => x"484a66c4",
  2377 => x"06a8b7c0",
  2378 => x"6e87d0c0",
  2379 => x"c480cc48",
  2380 => x"8ac158a6",
  2381 => x"01aab7c0",
  2382 => x"6e87f0ff",
  2383 => x"c24bbf97",
  2384 => x"d1c0028b",
  2385 => x"c0058b87",
  2386 => x"4a6e87d7",
  2387 => x"496a82c8",
  2388 => x"c087c2f5",
  2389 => x"4b6e87cb",
  2390 => x"4b6b83c8",
  2391 => x"734966c4",
  2392 => x"029d750f",
  2393 => x"6d87e9c0",
  2394 => x"87e4c002",
  2395 => x"dbff496d",
  2396 => x"497087ed",
  2397 => x"c00299c1",
  2398 => x"a5c487cb",
  2399 => x"ceecc24b",
  2400 => x"4b6b49bf",
  2401 => x"0285c80f",
  2402 => x"6d87c5c0",
  2403 => x"87dcff05",
  2404 => x"c00266c8",
  2405 => x"ecc287c8",
  2406 => x"f149bfce",
  2407 => x"8ef487e0",
  2408 => x"5887eaf3",
  2409 => x"1d141112",
  2410 => x"5a231c1b",
  2411 => x"f5949159",
  2412 => x"00f4ebf2",
  2413 => x"00000000",
  2414 => x"00000000",
  2415 => x"58000000",
  2416 => x"1d111412",
  2417 => x"5a231c1b",
  2418 => x"f5919459",
  2419 => x"00f4ebf2",
  2420 => x"000025d4",
  2421 => x"4f545541",
  2422 => x"544f4f42",
  2423 => x"0053454e",
  2424 => x"000019d4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
