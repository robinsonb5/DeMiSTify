library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dce7c287",
    12 => x"48c0c44e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90588",
    17 => x"49dce7c2",
    18 => x"48ecd2c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"ead2c287",
    25 => x"e6d2c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e0c187f7",
    29 => x"d2c287d9",
    30 => x"d2c24dea",
    31 => x"ad744cea",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"c04b710e",
    37 => x"9a4a134c",
    38 => x"7287cd02",
    39 => x"87e0c049",
    40 => x"4a1384c1",
    41 => x"87f3059a",
    42 => x"4c264874",
    43 => x"4f264b26",
    44 => x"8148731e",
    45 => x"c502a973",
    46 => x"05531287",
    47 => x"4f2687f6",
    48 => x"c0ff1e1e",
    49 => x"c4486a4a",
    50 => x"a6c498c0",
    51 => x"02987058",
    52 => x"7a7187f3",
    53 => x"4f262648",
    54 => x"ff1e731e",
    55 => x"ffc34bd4",
    56 => x"c34a6b7b",
    57 => x"496b7bff",
    58 => x"b17232c8",
    59 => x"6b7bffc3",
    60 => x"7131c84a",
    61 => x"7bffc3b2",
    62 => x"32c8496b",
    63 => x"4871b172",
    64 => x"4d2687c4",
    65 => x"4b264c26",
    66 => x"5e0e4f26",
    67 => x"0e5d5c5b",
    68 => x"d4ff4a71",
    69 => x"c348724c",
    70 => x"7c7098ff",
    71 => x"bfecd2c2",
    72 => x"d087c805",
    73 => x"30c94866",
    74 => x"d058a6d4",
    75 => x"29d84966",
    76 => x"ffc34871",
    77 => x"d07c7098",
    78 => x"29d04966",
    79 => x"ffc34871",
    80 => x"d07c7098",
    81 => x"29c84966",
    82 => x"ffc34871",
    83 => x"d07c7098",
    84 => x"ffc34866",
    85 => x"727c7098",
    86 => x"7129d049",
    87 => x"98ffc348",
    88 => x"4b6c7c70",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87fffd",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487dffd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c1fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87defc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"49e3c878",
   125 => x"d387d5fa",
   126 => x"c01ec04b",
   127 => x"c1c1f0ff",
   128 => x"87c6fc49",
   129 => x"987086c4",
   130 => x"ff87ca05",
   131 => x"ffc348d4",
   132 => x"cb48c178",
   133 => x"87ebfd87",
   134 => x"ff058bc1",
   135 => x"48c087db",
   136 => x"4387e3fb",
   137 => x"5300444d",
   138 => x"20434844",
   139 => x"6c696166",
   140 => x"49000a21",
   141 => x"00525245",
   142 => x"00495053",
   143 => x"74697257",
   144 => x"61662065",
   145 => x"64656c69",
   146 => x"5e0e000a",
   147 => x"ff0e5c5b",
   148 => x"eefc4cd4",
   149 => x"1eeac687",
   150 => x"c1f0e1c0",
   151 => x"e9fa49c8",
   152 => x"c186c487",
   153 => x"87c802a8",
   154 => x"c087fdfd",
   155 => x"87e8c148",
   156 => x"7087e5f9",
   157 => x"ffffcf49",
   158 => x"a9eac699",
   159 => x"fd87c802",
   160 => x"48c087e6",
   161 => x"c387d1c1",
   162 => x"f1c07cff",
   163 => x"87c7fc4b",
   164 => x"c0029870",
   165 => x"1ec087eb",
   166 => x"c1f0ffc0",
   167 => x"e9f949fa",
   168 => x"7086c487",
   169 => x"87d90598",
   170 => x"6c7cffc3",
   171 => x"7cffc349",
   172 => x"c17c7c7c",
   173 => x"c40299c0",
   174 => x"db48c187",
   175 => x"d748c087",
   176 => x"05abc287",
   177 => x"e7c887ca",
   178 => x"87c0f749",
   179 => x"87c848c0",
   180 => x"fe058bc1",
   181 => x"48c087f7",
   182 => x"0e87e9f8",
   183 => x"5d5c5b5e",
   184 => x"d0ff1e0e",
   185 => x"c0c0c84d",
   186 => x"ecd2c24b",
   187 => x"c878c148",
   188 => x"d7f649f8",
   189 => x"6d4cc787",
   190 => x"c4987348",
   191 => x"987058a6",
   192 => x"6d87cc02",
   193 => x"c4987348",
   194 => x"987058a6",
   195 => x"c287f405",
   196 => x"87eff97d",
   197 => x"9873486d",
   198 => x"7058a6c4",
   199 => x"87cc0298",
   200 => x"9873486d",
   201 => x"7058a6c4",
   202 => x"87f40598",
   203 => x"1ec07dc3",
   204 => x"c1d0e5c0",
   205 => x"d1f749c0",
   206 => x"c186c487",
   207 => x"87c105a8",
   208 => x"05acc24c",
   209 => x"f3c887cb",
   210 => x"87c0f549",
   211 => x"cec148c0",
   212 => x"058cc187",
   213 => x"fb87e0fe",
   214 => x"d2c287f0",
   215 => x"987058f0",
   216 => x"c187cd05",
   217 => x"f0ffc01e",
   218 => x"f649d0c1",
   219 => x"86c487dc",
   220 => x"c348d4ff",
   221 => x"ddc578ff",
   222 => x"f4d2c287",
   223 => x"73486d58",
   224 => x"58a6c498",
   225 => x"cc029870",
   226 => x"73486d87",
   227 => x"58a6c498",
   228 => x"f4059870",
   229 => x"ff7dc287",
   230 => x"ffc348d4",
   231 => x"2648c178",
   232 => x"0e87dff5",
   233 => x"5d5c5b5e",
   234 => x"c0c81e0e",
   235 => x"4cc04bc0",
   236 => x"dfcdeec5",
   237 => x"5ca6c44a",
   238 => x"c34cd4ff",
   239 => x"486c7cff",
   240 => x"05a8fec3",
   241 => x"7187c0c2",
   242 => x"e2c00599",
   243 => x"bfd0ff87",
   244 => x"c4987348",
   245 => x"987058a6",
   246 => x"ff87ce02",
   247 => x"7348bfd0",
   248 => x"58a6c498",
   249 => x"f2059870",
   250 => x"48d0ff87",
   251 => x"d478d1c4",
   252 => x"b7c04866",
   253 => x"e0c006a8",
   254 => x"7cffc387",
   255 => x"99714a6c",
   256 => x"7187c702",
   257 => x"0a7a970a",
   258 => x"66d481c1",
   259 => x"d888c148",
   260 => x"b7c058a6",
   261 => x"e0ff01a8",
   262 => x"7cffc387",
   263 => x"0599717c",
   264 => x"ff87e1c0",
   265 => x"7348bfd0",
   266 => x"58a6c498",
   267 => x"ce029870",
   268 => x"bfd0ff87",
   269 => x"c4987348",
   270 => x"987058a6",
   271 => x"ff87f205",
   272 => x"78d048d0",
   273 => x"c17e4ac1",
   274 => x"eefd058a",
   275 => x"26486e87",
   276 => x"0e87eff2",
   277 => x"0e5c5b5e",
   278 => x"c84a711e",
   279 => x"c04bc0c0",
   280 => x"48d4ff4c",
   281 => x"ff78ffc3",
   282 => x"7348bfd0",
   283 => x"58a6c498",
   284 => x"ce029870",
   285 => x"bfd0ff87",
   286 => x"c4987348",
   287 => x"987058a6",
   288 => x"ff87f205",
   289 => x"c3c448d0",
   290 => x"48d4ff78",
   291 => x"7278ffc3",
   292 => x"f0ffc01e",
   293 => x"f149d1c1",
   294 => x"86c487f0",
   295 => x"c0059870",
   296 => x"c0c887ee",
   297 => x"4966d41e",
   298 => x"c487f8fb",
   299 => x"ff4c7086",
   300 => x"7348bfd0",
   301 => x"58a6c498",
   302 => x"ce029870",
   303 => x"bfd0ff87",
   304 => x"c4987348",
   305 => x"987058a6",
   306 => x"ff87f205",
   307 => x"78c248d0",
   308 => x"f0264874",
   309 => x"5e0e87ee",
   310 => x"0e5d5c5b",
   311 => x"ffc01ec0",
   312 => x"49c9c1f0",
   313 => x"d287e3f0",
   314 => x"fad2c21e",
   315 => x"87f3fa49",
   316 => x"4cc086c8",
   317 => x"b7d284c1",
   318 => x"87f804ac",
   319 => x"97fad2c2",
   320 => x"c0c349bf",
   321 => x"a9c0c199",
   322 => x"87e7c005",
   323 => x"97c1d3c2",
   324 => x"31d049bf",
   325 => x"97c2d3c2",
   326 => x"32c84abf",
   327 => x"d3c2b172",
   328 => x"4abf97c3",
   329 => x"cf4c71b1",
   330 => x"9cffffff",
   331 => x"34ca84c1",
   332 => x"c287e7c1",
   333 => x"bf97c3d3",
   334 => x"c631c149",
   335 => x"c4d3c299",
   336 => x"c74abf97",
   337 => x"b1722ab7",
   338 => x"97ffd2c2",
   339 => x"cf4d4abf",
   340 => x"c0d3c29d",
   341 => x"c34abf97",
   342 => x"c232ca9a",
   343 => x"bf97c1d3",
   344 => x"7333c24b",
   345 => x"c2d3c2b2",
   346 => x"c34bbf97",
   347 => x"b7c69bc0",
   348 => x"c2b2732b",
   349 => x"7148c181",
   350 => x"c1497030",
   351 => x"70307548",
   352 => x"c14c724d",
   353 => x"c8947184",
   354 => x"06adb7c0",
   355 => x"34c187cc",
   356 => x"c0c82db7",
   357 => x"ff01adb7",
   358 => x"487487f4",
   359 => x"0e87e3ed",
   360 => x"0e5c5b5e",
   361 => x"4cc04b71",
   362 => x"c04866d0",
   363 => x"c006a8b7",
   364 => x"4a1387e3",
   365 => x"bf9766cc",
   366 => x"4866cc49",
   367 => x"a6d080c1",
   368 => x"aab77158",
   369 => x"c187c402",
   370 => x"c187cc48",
   371 => x"b766d084",
   372 => x"ddff04ac",
   373 => x"c248c087",
   374 => x"264d2687",
   375 => x"264b264c",
   376 => x"5b5e0e4f",
   377 => x"c20e5d5c",
   378 => x"c048e0db",
   379 => x"d8d3c278",
   380 => x"f949c01e",
   381 => x"86c487dd",
   382 => x"c5059870",
   383 => x"c848c087",
   384 => x"4bc087ef",
   385 => x"48d8e0c2",
   386 => x"1ec878c1",
   387 => x"1efde0c0",
   388 => x"49ced4c2",
   389 => x"c887c8fe",
   390 => x"05987086",
   391 => x"e0c287c6",
   392 => x"78c048d8",
   393 => x"e1c01ec8",
   394 => x"d4c21ec6",
   395 => x"eefd49ea",
   396 => x"7086c887",
   397 => x"87c60598",
   398 => x"48d8e0c2",
   399 => x"e0c278c0",
   400 => x"c002bfd8",
   401 => x"dac287fa",
   402 => x"c24bbfde",
   403 => x"bf9fd6db",
   404 => x"ead6c54a",
   405 => x"87c705aa",
   406 => x"bfdedac2",
   407 => x"ca87cc4b",
   408 => x"02aad5e9",
   409 => x"48c087c5",
   410 => x"c287c6c7",
   411 => x"731ed8d3",
   412 => x"87dff749",
   413 => x"987086c4",
   414 => x"c087c505",
   415 => x"87f1c648",
   416 => x"e1c01ec8",
   417 => x"d4c21ecf",
   418 => x"d2fc49ea",
   419 => x"7086c887",
   420 => x"87c80598",
   421 => x"48e0dbc2",
   422 => x"87da78c1",
   423 => x"e1c01ec8",
   424 => x"d4c21ed8",
   425 => x"f6fb49ce",
   426 => x"7086c887",
   427 => x"c5c00298",
   428 => x"c548c087",
   429 => x"dbc287fb",
   430 => x"49bf97d6",
   431 => x"05a9d5c1",
   432 => x"c287cdc0",
   433 => x"bf97d7db",
   434 => x"a9eac249",
   435 => x"87c5c002",
   436 => x"dcc548c0",
   437 => x"d8d3c287",
   438 => x"c34cbf97",
   439 => x"c002ace9",
   440 => x"ebc387cc",
   441 => x"c5c002ac",
   442 => x"c548c087",
   443 => x"d3c287c3",
   444 => x"49bf97e3",
   445 => x"ccc00599",
   446 => x"e4d3c287",
   447 => x"c249bf97",
   448 => x"c5c002a9",
   449 => x"c448c087",
   450 => x"d3c287e7",
   451 => x"48bf97e5",
   452 => x"58dcdbc2",
   453 => x"dbc288c1",
   454 => x"d3c258e0",
   455 => x"49bf97e6",
   456 => x"d3c28173",
   457 => x"4abf97e7",
   458 => x"7135c84d",
   459 => x"f8dfc285",
   460 => x"e8d3c25d",
   461 => x"c248bf97",
   462 => x"c258cce0",
   463 => x"02bfe0db",
   464 => x"c887dcc2",
   465 => x"f4e0c01e",
   466 => x"ead4c21e",
   467 => x"87cff949",
   468 => x"987086c8",
   469 => x"87c5c002",
   470 => x"d4c348c0",
   471 => x"d8dbc287",
   472 => x"c4484abf",
   473 => x"e8dbc230",
   474 => x"c8e0c258",
   475 => x"fdd3c25a",
   476 => x"c849bf97",
   477 => x"fcd3c231",
   478 => x"a14bbf97",
   479 => x"fed3c249",
   480 => x"d04bbf97",
   481 => x"49a17333",
   482 => x"97ffd3c2",
   483 => x"33d84bbf",
   484 => x"c249a173",
   485 => x"c259d0e0",
   486 => x"91bfc8e0",
   487 => x"bff4dfc2",
   488 => x"fcdfc281",
   489 => x"c5d4c259",
   490 => x"c84bbf97",
   491 => x"c4d4c233",
   492 => x"a34cbf97",
   493 => x"c6d4c24b",
   494 => x"d04cbf97",
   495 => x"4ba37434",
   496 => x"97c7d4c2",
   497 => x"9ccf4cbf",
   498 => x"a37434d8",
   499 => x"c0e0c24b",
   500 => x"738bc25b",
   501 => x"c0e0c292",
   502 => x"78a17248",
   503 => x"c287cbc1",
   504 => x"bf97ead3",
   505 => x"c231c849",
   506 => x"bf97e9d3",
   507 => x"c249a14a",
   508 => x"c559e8db",
   509 => x"81ffc731",
   510 => x"e0c229c9",
   511 => x"d3c259c8",
   512 => x"4abf97ef",
   513 => x"d3c232c8",
   514 => x"4bbf97ee",
   515 => x"e0c24aa2",
   516 => x"e0c25ad0",
   517 => x"7592bfc8",
   518 => x"c4e0c282",
   519 => x"fcdfc25a",
   520 => x"c278c048",
   521 => x"7248f8df",
   522 => x"49c078a1",
   523 => x"c187f7c7",
   524 => x"87e5f648",
   525 => x"33544146",
   526 => x"20202032",
   527 => x"54414600",
   528 => x"20203631",
   529 => x"41460020",
   530 => x"20323354",
   531 => x"46002020",
   532 => x"32335441",
   533 => x"00202020",
   534 => x"31544146",
   535 => x"20202036",
   536 => x"5b5e0e00",
   537 => x"710e5d5c",
   538 => x"e0dbc24a",
   539 => x"87cc02bf",
   540 => x"b7c74b72",
   541 => x"c14d722b",
   542 => x"87ca9dff",
   543 => x"b7c84b72",
   544 => x"c34d722b",
   545 => x"d3c29dff",
   546 => x"dfc21ed8",
   547 => x"7349bff4",
   548 => x"feee7181",
   549 => x"7086c487",
   550 => x"87c50598",
   551 => x"e6c048c0",
   552 => x"e0dbc287",
   553 => x"87d202bf",
   554 => x"91c44975",
   555 => x"81d8d3c2",
   556 => x"ffcf4c69",
   557 => x"9cffffff",
   558 => x"497587cb",
   559 => x"d3c291c2",
   560 => x"699f81d8",
   561 => x"f448744c",
   562 => x"5e0e87cf",
   563 => x"0e5d5c5b",
   564 => x"4c7186f4",
   565 => x"e0c24bc0",
   566 => x"c47ebfd0",
   567 => x"e0c248a6",
   568 => x"c878bfd4",
   569 => x"78c048a6",
   570 => x"bfe4dbc2",
   571 => x"06a8c048",
   572 => x"c887ddc2",
   573 => x"99cf4966",
   574 => x"c287d805",
   575 => x"c81ed8d3",
   576 => x"c1484966",
   577 => x"58a6cc80",
   578 => x"c487c8ed",
   579 => x"d8d3c286",
   580 => x"c087c34b",
   581 => x"6b9783e0",
   582 => x"c1029a4a",
   583 => x"e5c387e1",
   584 => x"dac102aa",
   585 => x"49a3cb87",
   586 => x"d8496997",
   587 => x"cec10599",
   588 => x"c01ecb87",
   589 => x"731e66e0",
   590 => x"87e3f149",
   591 => x"987086c8",
   592 => x"87fbc005",
   593 => x"c44aa3dc",
   594 => x"796a49a4",
   595 => x"c849a3da",
   596 => x"699f4da4",
   597 => x"dbc27d48",
   598 => x"d302bfe0",
   599 => x"49a3d487",
   600 => x"c049699f",
   601 => x"7199ffff",
   602 => x"c430d048",
   603 => x"87c258a6",
   604 => x"486e7ec0",
   605 => x"7d70806d",
   606 => x"48c17cc0",
   607 => x"c887c5c1",
   608 => x"80c14866",
   609 => x"c258a6cc",
   610 => x"a8bfe4db",
   611 => x"87e3fd04",
   612 => x"bfe0dbc2",
   613 => x"87eac002",
   614 => x"c4fb496e",
   615 => x"58a6c487",
   616 => x"ffcf4970",
   617 => x"99f8ffff",
   618 => x"87d602a9",
   619 => x"89c24970",
   620 => x"bfd8dbc2",
   621 => x"f8dfc291",
   622 => x"807148bf",
   623 => x"fc58a6c8",
   624 => x"48c087e1",
   625 => x"d0f08ef4",
   626 => x"1e731e87",
   627 => x"496a4a71",
   628 => x"7a7181c1",
   629 => x"bfdcdbc2",
   630 => x"87cb0599",
   631 => x"6b4ba2c8",
   632 => x"87fdf949",
   633 => x"c17b4970",
   634 => x"87f1ef48",
   635 => x"711e731e",
   636 => x"f8dfc24b",
   637 => x"a3c849bf",
   638 => x"c24a6a4a",
   639 => x"d8dbc28a",
   640 => x"a17292bf",
   641 => x"dcdbc249",
   642 => x"9a6b4abf",
   643 => x"c849a172",
   644 => x"e8711e66",
   645 => x"86c487fd",
   646 => x"c4059870",
   647 => x"c248c087",
   648 => x"ee48c187",
   649 => x"5e0e87f7",
   650 => x"710e5c5b",
   651 => x"724bc04a",
   652 => x"e0c0029a",
   653 => x"49a2da87",
   654 => x"c24b699f",
   655 => x"02bfe0db",
   656 => x"a2d487cf",
   657 => x"49699f49",
   658 => x"ffffc04c",
   659 => x"c234d09c",
   660 => x"744cc087",
   661 => x"029b73b3",
   662 => x"c24a87df",
   663 => x"d8dbc28a",
   664 => x"c29249bf",
   665 => x"48bff8df",
   666 => x"e0c28072",
   667 => x"487158d8",
   668 => x"dbc230c4",
   669 => x"e9c058e8",
   670 => x"fcdfc287",
   671 => x"e0c24bbf",
   672 => x"e0c248d4",
   673 => x"c278bfc0",
   674 => x"02bfe0db",
   675 => x"dbc287c9",
   676 => x"c449bfd8",
   677 => x"c287c731",
   678 => x"49bfc4e0",
   679 => x"dbc231c4",
   680 => x"e0c259e8",
   681 => x"f2ec5bd4",
   682 => x"5b5e0e87",
   683 => x"f40e5d5c",
   684 => x"9a4a7186",
   685 => x"c287de02",
   686 => x"c048d4d3",
   687 => x"ccd3c278",
   688 => x"d4e0c248",
   689 => x"d3c278bf",
   690 => x"e0c248d0",
   691 => x"c078bfd0",
   692 => x"c048fff1",
   693 => x"e4dbc278",
   694 => x"d3c249bf",
   695 => x"714abfd4",
   696 => x"cbc403aa",
   697 => x"cf497287",
   698 => x"e0c00599",
   699 => x"d8d3c287",
   700 => x"ccd3c21e",
   701 => x"d3c249bf",
   702 => x"a1c148cc",
   703 => x"d2e57178",
   704 => x"c086c487",
   705 => x"c248fbf1",
   706 => x"cc78d8d3",
   707 => x"fbf1c087",
   708 => x"e0c048bf",
   709 => x"fff1c080",
   710 => x"d4d3c258",
   711 => x"80c148bf",
   712 => x"58d8d3c2",
   713 => x"000c7b27",
   714 => x"bf97bf00",
   715 => x"c2029c4c",
   716 => x"e5c387ee",
   717 => x"e7c202ac",
   718 => x"fbf1c087",
   719 => x"a3cb4bbf",
   720 => x"cf4d1149",
   721 => x"d6c105ad",
   722 => x"df497487",
   723 => x"cd89c199",
   724 => x"e8dbc291",
   725 => x"4aa3c181",
   726 => x"a3c35112",
   727 => x"c551124a",
   728 => x"51124aa3",
   729 => x"124aa3c7",
   730 => x"4aa3c951",
   731 => x"a3ce5112",
   732 => x"d051124a",
   733 => x"51124aa3",
   734 => x"124aa3d2",
   735 => x"4aa3d451",
   736 => x"a3d65112",
   737 => x"d851124a",
   738 => x"51124aa3",
   739 => x"124aa3dc",
   740 => x"4aa3de51",
   741 => x"f1c05112",
   742 => x"78c148ff",
   743 => x"7587c1c1",
   744 => x"0599c849",
   745 => x"7587f3c0",
   746 => x"0599d049",
   747 => x"66dc87d0",
   748 => x"87cac002",
   749 => x"66dc4973",
   750 => x"0298700f",
   751 => x"f1c087dc",
   752 => x"c005bfff",
   753 => x"dbc287c6",
   754 => x"50c048e8",
   755 => x"48fff1c0",
   756 => x"f1c078c0",
   757 => x"c248bffb",
   758 => x"f1c087dc",
   759 => x"78c048ff",
   760 => x"bfe4dbc2",
   761 => x"d4d3c249",
   762 => x"aa714abf",
   763 => x"87f5fb04",
   764 => x"bfd4e0c2",
   765 => x"87c8c005",
   766 => x"bfe0dbc2",
   767 => x"87f4c102",
   768 => x"bfd0d3c2",
   769 => x"87d9f149",
   770 => x"58d4d3c2",
   771 => x"dbc27e70",
   772 => x"c002bfe0",
   773 => x"496e87dd",
   774 => x"ffffffcf",
   775 => x"02a999f8",
   776 => x"c487c8c0",
   777 => x"78c048a6",
   778 => x"c487e6c0",
   779 => x"78c148a6",
   780 => x"6e87dec0",
   781 => x"f8ffcf49",
   782 => x"c002a999",
   783 => x"a6c887c8",
   784 => x"c078c048",
   785 => x"a6c887c5",
   786 => x"c478c148",
   787 => x"66c848a6",
   788 => x"0566c478",
   789 => x"6e87ddc0",
   790 => x"c289c249",
   791 => x"91bfd8db",
   792 => x"bff8dfc2",
   793 => x"c2807148",
   794 => x"c258d0d3",
   795 => x"c048d4d3",
   796 => x"87e1f978",
   797 => x"8ef448c0",
   798 => x"0087dee5",
   799 => x"00000000",
   800 => x"1e000000",
   801 => x"c348d4ff",
   802 => x"496878ff",
   803 => x"87c60299",
   804 => x"05a9fbc0",
   805 => x"487187ee",
   806 => x"5e0e4f26",
   807 => x"710e5c5b",
   808 => x"ff4bc04a",
   809 => x"ffc348d4",
   810 => x"99496878",
   811 => x"87c1c102",
   812 => x"02a9ecc0",
   813 => x"c087fac0",
   814 => x"c002a9fb",
   815 => x"66cc87f3",
   816 => x"cc03abb7",
   817 => x"0266d087",
   818 => x"097287c7",
   819 => x"c1097997",
   820 => x"02997182",
   821 => x"83c187c2",
   822 => x"c348d4ff",
   823 => x"496878ff",
   824 => x"87cd0299",
   825 => x"02a9ecc0",
   826 => x"fbc087c7",
   827 => x"cdff05a9",
   828 => x"0266d087",
   829 => x"97c087c3",
   830 => x"a9fbc07a",
   831 => x"7387c705",
   832 => x"8c0cc04c",
   833 => x"4c7387c2",
   834 => x"87c24874",
   835 => x"4c264d26",
   836 => x"4f264b26",
   837 => x"48d4ff1e",
   838 => x"6878ffc3",
   839 => x"b7f0c049",
   840 => x"87ca04a9",
   841 => x"a9b7f9c0",
   842 => x"c087c301",
   843 => x"c1c189f0",
   844 => x"ca04a9b7",
   845 => x"b7c6c187",
   846 => x"87c301a9",
   847 => x"7189f7c0",
   848 => x"0e4f2648",
   849 => x"5d5c5b5e",
   850 => x"7186f40e",
   851 => x"4bd4ff4c",
   852 => x"c37e4dc0",
   853 => x"d0ff7bff",
   854 => x"c0c848bf",
   855 => x"a6c898c0",
   856 => x"02987058",
   857 => x"d0ff87d0",
   858 => x"c0c848bf",
   859 => x"a6c898c0",
   860 => x"05987058",
   861 => x"d0ff87f0",
   862 => x"78e1c048",
   863 => x"c2fc7bd4",
   864 => x"99497087",
   865 => x"87c7c102",
   866 => x"c87bffc3",
   867 => x"786b48a6",
   868 => x"c04866c8",
   869 => x"c802a8fb",
   870 => x"f0e0c287",
   871 => x"eec002bf",
   872 => x"714dc187",
   873 => x"e6c00299",
   874 => x"a9fbc087",
   875 => x"fb87c302",
   876 => x"ffc387d1",
   877 => x"c1496b7b",
   878 => x"cc05a9c6",
   879 => x"7bffc387",
   880 => x"48a6c87b",
   881 => x"49c0786b",
   882 => x"0599714d",
   883 => x"7587daff",
   884 => x"dec1059d",
   885 => x"7bffc387",
   886 => x"ffc34a6b",
   887 => x"48a6c47b",
   888 => x"486e786b",
   889 => x"a6c480c1",
   890 => x"49a4c858",
   891 => x"c8496997",
   892 => x"da05a966",
   893 => x"49a4c987",
   894 => x"aa496997",
   895 => x"ca87d005",
   896 => x"699749a4",
   897 => x"a966c449",
   898 => x"c187c405",
   899 => x"c887d64d",
   900 => x"ecc04866",
   901 => x"87c902a8",
   902 => x"c04866c8",
   903 => x"c405a8fb",
   904 => x"c17ec087",
   905 => x"7bffc34d",
   906 => x"6b48a6c8",
   907 => x"029d7578",
   908 => x"ff87e2fe",
   909 => x"c848bfd0",
   910 => x"c898c0c0",
   911 => x"987058a6",
   912 => x"ff87d002",
   913 => x"c848bfd0",
   914 => x"c898c0c0",
   915 => x"987058a6",
   916 => x"ff87f005",
   917 => x"e0c048d0",
   918 => x"f4486e78",
   919 => x"87ecfa8e",
   920 => x"5c5b5e0e",
   921 => x"86f40e5d",
   922 => x"ff59a6c4",
   923 => x"c0c84cd0",
   924 => x"1e6e4bc0",
   925 => x"49f4e0c2",
   926 => x"c487cfe9",
   927 => x"02987086",
   928 => x"c287f7c5",
   929 => x"4dbff8e0",
   930 => x"f6fa496e",
   931 => x"58a6c887",
   932 => x"9873486c",
   933 => x"7058a6cc",
   934 => x"87cc0298",
   935 => x"9873486c",
   936 => x"7058a6c4",
   937 => x"87f40598",
   938 => x"d4ff7cc5",
   939 => x"78d5c148",
   940 => x"bff0e0c2",
   941 => x"c481c149",
   942 => x"8ac14a66",
   943 => x"487232c6",
   944 => x"d4ffb071",
   945 => x"486c7808",
   946 => x"a6c49873",
   947 => x"02987058",
   948 => x"486c87cc",
   949 => x"a6c49873",
   950 => x"05987058",
   951 => x"7cc487f4",
   952 => x"c348d4ff",
   953 => x"486c78ff",
   954 => x"a6c49873",
   955 => x"02987058",
   956 => x"486c87cc",
   957 => x"a6c49873",
   958 => x"05987058",
   959 => x"7cc587f4",
   960 => x"c148d4ff",
   961 => x"78c178d3",
   962 => x"9873486c",
   963 => x"7058a6c4",
   964 => x"87cc0298",
   965 => x"9873486c",
   966 => x"7058a6c4",
   967 => x"87f40598",
   968 => x"9d757cc4",
   969 => x"87d0c202",
   970 => x"7ed8d3c2",
   971 => x"f4e0c21e",
   972 => x"87f8ea49",
   973 => x"987086c4",
   974 => x"c087c505",
   975 => x"87fcc248",
   976 => x"adb7c0c8",
   977 => x"4a87c404",
   978 => x"7587c48d",
   979 => x"6c4dc04a",
   980 => x"c8987348",
   981 => x"987058a6",
   982 => x"6c87cc02",
   983 => x"c8987348",
   984 => x"987058a6",
   985 => x"cd87f405",
   986 => x"48d4ff7c",
   987 => x"7278d4c1",
   988 => x"718ac149",
   989 => x"87d90299",
   990 => x"48bf976e",
   991 => x"7808d4ff",
   992 => x"80c1486e",
   993 => x"7258a6c4",
   994 => x"718ac149",
   995 => x"e7ff0599",
   996 => x"73486c87",
   997 => x"58a6c498",
   998 => x"cc029870",
   999 => x"73486c87",
  1000 => x"58a6c498",
  1001 => x"f4059870",
  1002 => x"c27cc487",
  1003 => x"e849f4e0",
  1004 => x"9d7587d7",
  1005 => x"87f0fd05",
  1006 => x"9873486c",
  1007 => x"7058a6c4",
  1008 => x"87cd0298",
  1009 => x"9873486c",
  1010 => x"7058a6c4",
  1011 => x"f3ff0598",
  1012 => x"ff7cc587",
  1013 => x"d3c148d4",
  1014 => x"6c78c078",
  1015 => x"c4987348",
  1016 => x"987058a6",
  1017 => x"6c87cd02",
  1018 => x"c4987348",
  1019 => x"987058a6",
  1020 => x"87f3ff05",
  1021 => x"48c17cc4",
  1022 => x"48c087c2",
  1023 => x"cbf48ef4",
  1024 => x"5b5e0e87",
  1025 => x"1e0e5d5c",
  1026 => x"4cc04b71",
  1027 => x"04abb74d",
  1028 => x"c087e9c0",
  1029 => x"751ec3f5",
  1030 => x"87c4029d",
  1031 => x"87c24ac0",
  1032 => x"49724ac1",
  1033 => x"c487c2ea",
  1034 => x"c158a686",
  1035 => x"c2056e84",
  1036 => x"c14c7387",
  1037 => x"acb77385",
  1038 => x"87d7ff06",
  1039 => x"f326486e",
  1040 => x"5e0e87ca",
  1041 => x"0e5d5c5b",
  1042 => x"494c711e",
  1043 => x"bfc4e1c2",
  1044 => x"87edfe81",
  1045 => x"029d4d70",
  1046 => x"c287fcc0",
  1047 => x"754be8db",
  1048 => x"ff49cb4a",
  1049 => x"7487c9c1",
  1050 => x"c291de49",
  1051 => x"7148d8e1",
  1052 => x"58a6c480",
  1053 => x"48e7c2c1",
  1054 => x"a1c8496e",
  1055 => x"7141204a",
  1056 => x"87f905aa",
  1057 => x"51105110",
  1058 => x"49745110",
  1059 => x"87fdc4c1",
  1060 => x"49e8dbc2",
  1061 => x"c187c9f7",
  1062 => x"c149f8e3",
  1063 => x"c187c0c6",
  1064 => x"2687cfc6",
  1065 => x"4c87e5f1",
  1066 => x"6964616f",
  1067 => x"2e2e676e",
  1068 => x"2080002e",
  1069 => x"6b636142",
  1070 => x"616f4c00",
  1071 => x"2e2a2064",
  1072 => x"203a0020",
  1073 => x"42208000",
  1074 => x"006b6361",
  1075 => x"78452080",
  1076 => x"53007469",
  1077 => x"6e492044",
  1078 => x"2e2e7469",
  1079 => x"004b4f00",
  1080 => x"544f4f42",
  1081 => x"20202020",
  1082 => x"004d4f52",
  1083 => x"711e731e",
  1084 => x"e1c2494b",
  1085 => x"fc81bfc4",
  1086 => x"4a7087c7",
  1087 => x"87c4029a",
  1088 => x"87e2e449",
  1089 => x"48c4e1c2",
  1090 => x"497378c0",
  1091 => x"ef87e9c1",
  1092 => x"731e87fe",
  1093 => x"c44b711e",
  1094 => x"c1024aa3",
  1095 => x"8ac187c8",
  1096 => x"8a87dc02",
  1097 => x"87f1c002",
  1098 => x"c4c1058a",
  1099 => x"c4e1c287",
  1100 => x"fcc002bf",
  1101 => x"88c14887",
  1102 => x"58c8e1c2",
  1103 => x"c287f2c0",
  1104 => x"49bfc4e1",
  1105 => x"e1c289d0",
  1106 => x"b7c059c8",
  1107 => x"e0c003a9",
  1108 => x"c4e1c287",
  1109 => x"d878c048",
  1110 => x"c4e1c287",
  1111 => x"80c148bf",
  1112 => x"58c8e1c2",
  1113 => x"e1c287cb",
  1114 => x"d048bfc4",
  1115 => x"c8e1c280",
  1116 => x"c3497358",
  1117 => x"87d8ee87",
  1118 => x"5c5b5e0e",
  1119 => x"86f00e5d",
  1120 => x"c259a6d0",
  1121 => x"c04dd8d3",
  1122 => x"48a6c44c",
  1123 => x"e1c278c0",
  1124 => x"c048bfc4",
  1125 => x"c106a8b7",
  1126 => x"d3c287c1",
  1127 => x"029848d8",
  1128 => x"c087f8c0",
  1129 => x"c81ec3f5",
  1130 => x"87c70266",
  1131 => x"c048a6c4",
  1132 => x"c487c578",
  1133 => x"78c148a6",
  1134 => x"e34966c4",
  1135 => x"86c487eb",
  1136 => x"84c14d70",
  1137 => x"c14866c4",
  1138 => x"58a6c880",
  1139 => x"bfc4e1c2",
  1140 => x"c603acb7",
  1141 => x"059d7587",
  1142 => x"c087c8ff",
  1143 => x"029d754c",
  1144 => x"c087dec3",
  1145 => x"c81ec3f5",
  1146 => x"87c70266",
  1147 => x"c048a6cc",
  1148 => x"cc87c578",
  1149 => x"78c148a6",
  1150 => x"e24966cc",
  1151 => x"86c487eb",
  1152 => x"026e58a6",
  1153 => x"4987e6c2",
  1154 => x"699781cb",
  1155 => x"0299d049",
  1156 => x"c187d6c1",
  1157 => x"744aecc3",
  1158 => x"c191cb49",
  1159 => x"7281f8e3",
  1160 => x"c381c879",
  1161 => x"497451ff",
  1162 => x"e1c291de",
  1163 => x"85714dd8",
  1164 => x"7d97c1c2",
  1165 => x"c049a5c1",
  1166 => x"dbc251e0",
  1167 => x"02bf97e8",
  1168 => x"84c187d2",
  1169 => x"c24ba5c2",
  1170 => x"db4ae8db",
  1171 => x"dff9fe49",
  1172 => x"87d9c187",
  1173 => x"c049a5cd",
  1174 => x"c284c151",
  1175 => x"4a6e4ba5",
  1176 => x"f9fe49cb",
  1177 => x"c4c187ca",
  1178 => x"cb497487",
  1179 => x"f8e3c191",
  1180 => x"c2c1c181",
  1181 => x"e8dbc279",
  1182 => x"d802bf97",
  1183 => x"de497487",
  1184 => x"c284c191",
  1185 => x"714bd8e1",
  1186 => x"e8dbc283",
  1187 => x"fe49dd4a",
  1188 => x"d887ddf8",
  1189 => x"de4b7487",
  1190 => x"d8e1c293",
  1191 => x"49a3cb83",
  1192 => x"84c151c0",
  1193 => x"cb4a6e73",
  1194 => x"c3f8fe49",
  1195 => x"4866c487",
  1196 => x"a6c880c1",
  1197 => x"acb7c758",
  1198 => x"87c5c003",
  1199 => x"e2fc056e",
  1200 => x"acb7c787",
  1201 => x"87d3c003",
  1202 => x"91de4974",
  1203 => x"81d8e1c2",
  1204 => x"84c151c0",
  1205 => x"04acb7c7",
  1206 => x"c187edff",
  1207 => x"c048cde5",
  1208 => x"c5e5c150",
  1209 => x"d3ccc148",
  1210 => x"c9e5c178",
  1211 => x"f2c2c148",
  1212 => x"d0e5c178",
  1213 => x"d2c4c148",
  1214 => x"4966cc78",
  1215 => x"87cdfbc0",
  1216 => x"c7e88ef0",
  1217 => x"4a711e87",
  1218 => x"5af4e0c2",
  1219 => x"e7f94972",
  1220 => x"1e4f2687",
  1221 => x"cb494a71",
  1222 => x"f8e3c191",
  1223 => x"1181c881",
  1224 => x"f0e0c248",
  1225 => x"a2f0c058",
  1226 => x"d3f6fe49",
  1227 => x"d549c087",
  1228 => x"4f2687c0",
  1229 => x"5c5b5e0e",
  1230 => x"86f00e5d",
  1231 => x"cb494d71",
  1232 => x"f8e3c191",
  1233 => x"7ea1ca81",
  1234 => x"c248a6c4",
  1235 => x"78bfe8e0",
  1236 => x"4abf976e",
  1237 => x"724b66c4",
  1238 => x"4aa1c82b",
  1239 => x"a6cc4812",
  1240 => x"c19b7058",
  1241 => x"9781c983",
  1242 => x"abb74969",
  1243 => x"c087c204",
  1244 => x"bf976e4b",
  1245 => x"4966c84a",
  1246 => x"b9ff3172",
  1247 => x"739966c4",
  1248 => x"7134724c",
  1249 => x"ece0c2b4",
  1250 => x"48d4ff5c",
  1251 => x"ff78ffc3",
  1252 => x"c848bfd0",
  1253 => x"d098c0c0",
  1254 => x"987058a6",
  1255 => x"ff87d002",
  1256 => x"c848bfd0",
  1257 => x"c498c0c0",
  1258 => x"987058a6",
  1259 => x"ff87f005",
  1260 => x"e1c048d0",
  1261 => x"48d4ff78",
  1262 => x"0c7078de",
  1263 => x"48740c7c",
  1264 => x"ff28b7c8",
  1265 => x"747808d4",
  1266 => x"28b7d048",
  1267 => x"7808d4ff",
  1268 => x"b7d84874",
  1269 => x"08d4ff28",
  1270 => x"bfd0ff78",
  1271 => x"c0c0c848",
  1272 => x"58a6c498",
  1273 => x"d0029870",
  1274 => x"bfd0ff87",
  1275 => x"c0c0c848",
  1276 => x"58a6c498",
  1277 => x"f0059870",
  1278 => x"48d0ff87",
  1279 => x"c778e0c0",
  1280 => x"c11ec01e",
  1281 => x"c21ef8e3",
  1282 => x"49bfece0",
  1283 => x"7587e1c1",
  1284 => x"f8f6c049",
  1285 => x"e38ee487",
  1286 => x"731e87f2",
  1287 => x"494b711e",
  1288 => x"7387d1fc",
  1289 => x"87ccfc49",
  1290 => x"1e87e5e3",
  1291 => x"4b711e73",
  1292 => x"024aa3c2",
  1293 => x"8ac187d5",
  1294 => x"c287db05",
  1295 => x"02bfc0e1",
  1296 => x"c14887d4",
  1297 => x"c4e1c288",
  1298 => x"c287cb58",
  1299 => x"48bfc0e1",
  1300 => x"e1c280c1",
  1301 => x"1ec758c4",
  1302 => x"e3c11ec0",
  1303 => x"e0c21ef8",
  1304 => x"cb49bfec",
  1305 => x"c0497387",
  1306 => x"f487e2f5",
  1307 => x"87e0e28e",
  1308 => x"5c5b5e0e",
  1309 => x"d8ff0e5d",
  1310 => x"59a6dc86",
  1311 => x"c048a6c8",
  1312 => x"c080c478",
  1313 => x"80c44d78",
  1314 => x"bfc0e1c2",
  1315 => x"48d4ff78",
  1316 => x"ff78ffc3",
  1317 => x"c848bfd0",
  1318 => x"c498c0c0",
  1319 => x"987058a6",
  1320 => x"ff87d002",
  1321 => x"c848bfd0",
  1322 => x"c498c0c0",
  1323 => x"987058a6",
  1324 => x"ff87f005",
  1325 => x"e1c048d0",
  1326 => x"48d4ff78",
  1327 => x"dfff78d4",
  1328 => x"d4ff87c1",
  1329 => x"78ffc348",
  1330 => x"ff48a6d4",
  1331 => x"d478bfd4",
  1332 => x"fbc04866",
  1333 => x"d1c102a8",
  1334 => x"66f8c087",
  1335 => x"6a82c44a",
  1336 => x"c11e727e",
  1337 => x"c448f9c2",
  1338 => x"a1c84966",
  1339 => x"7141204a",
  1340 => x"87f905aa",
  1341 => x"4a265110",
  1342 => x"4866f8c0",
  1343 => x"78c5ccc1",
  1344 => x"81c7496a",
  1345 => x"c15166d4",
  1346 => x"6a1ed81e",
  1347 => x"ff81c849",
  1348 => x"c887c7de",
  1349 => x"4866d086",
  1350 => x"01a8b7c0",
  1351 => x"4dc187c4",
  1352 => x"66d087c8",
  1353 => x"d488c148",
  1354 => x"66d458a6",
  1355 => x"87e5ca02",
  1356 => x"b766c0c1",
  1357 => x"dcca03ad",
  1358 => x"48d4ff87",
  1359 => x"d478ffc3",
  1360 => x"d4ff48a6",
  1361 => x"66d478bf",
  1362 => x"88c6c148",
  1363 => x"7058a6c4",
  1364 => x"e6c00298",
  1365 => x"88c94887",
  1366 => x"7058a6c4",
  1367 => x"cdc40298",
  1368 => x"88c14887",
  1369 => x"7058a6c4",
  1370 => x"e0c10298",
  1371 => x"88c44887",
  1372 => x"987058a6",
  1373 => x"87f6c302",
  1374 => x"d887c4c9",
  1375 => x"c2c10566",
  1376 => x"48d4ff87",
  1377 => x"c078ffc3",
  1378 => x"751eca1e",
  1379 => x"c193cb4b",
  1380 => x"c48366c0",
  1381 => x"496c4ca3",
  1382 => x"87fedbff",
  1383 => x"1ede1ec1",
  1384 => x"dbff496c",
  1385 => x"86d087f4",
  1386 => x"7bc5ccc1",
  1387 => x"adb766d0",
  1388 => x"c187c504",
  1389 => x"87cec885",
  1390 => x"c14866d0",
  1391 => x"58a6d488",
  1392 => x"ff87c3c8",
  1393 => x"d887fcda",
  1394 => x"f9c758a6",
  1395 => x"c3ddff87",
  1396 => x"58a6cc87",
  1397 => x"a8b766cc",
  1398 => x"cc87c606",
  1399 => x"66c848a6",
  1400 => x"efdcff78",
  1401 => x"a8ecc087",
  1402 => x"87c2c205",
  1403 => x"c10566d8",
  1404 => x"497587f2",
  1405 => x"f8c091cb",
  1406 => x"a1c48166",
  1407 => x"c84c6a4a",
  1408 => x"66c84aa1",
  1409 => x"d3ccc152",
  1410 => x"48d4ff79",
  1411 => x"d478ffc3",
  1412 => x"d4ff48a6",
  1413 => x"66d478bf",
  1414 => x"87e8c002",
  1415 => x"a8fbc048",
  1416 => x"87e0c002",
  1417 => x"7c9766d4",
  1418 => x"d4ff84c1",
  1419 => x"78ffc348",
  1420 => x"ff48a6d4",
  1421 => x"d478bfd4",
  1422 => x"87c80266",
  1423 => x"a8fbc048",
  1424 => x"87e0ff05",
  1425 => x"c254e0c0",
  1426 => x"97c054c1",
  1427 => x"b766d07c",
  1428 => x"87c504ad",
  1429 => x"edc585c1",
  1430 => x"4866d087",
  1431 => x"a6d488c1",
  1432 => x"87e2c558",
  1433 => x"87dbd8ff",
  1434 => x"c558a6d8",
  1435 => x"66c887d8",
  1436 => x"a866d848",
  1437 => x"87fdc405",
  1438 => x"c048a6dc",
  1439 => x"d3daff78",
  1440 => x"58a6d887",
  1441 => x"87ccdaff",
  1442 => x"58a6e4c0",
  1443 => x"05a8ecc0",
  1444 => x"c087cac0",
  1445 => x"d448a6e0",
  1446 => x"c6c07866",
  1447 => x"48d4ff87",
  1448 => x"7578ffc3",
  1449 => x"c091cb49",
  1450 => x"714866f8",
  1451 => x"58a6c480",
  1452 => x"81ca496e",
  1453 => x"c05166d4",
  1454 => x"c14966e0",
  1455 => x"8966d481",
  1456 => x"307148c1",
  1457 => x"89c14970",
  1458 => x"82c84a6e",
  1459 => x"79970972",
  1460 => x"e8e0c209",
  1461 => x"66d449bf",
  1462 => x"6a9729b7",
  1463 => x"9871484a",
  1464 => x"58a6e8c0",
  1465 => x"80c4486e",
  1466 => x"c458a6c8",
  1467 => x"d84cbf66",
  1468 => x"66c84866",
  1469 => x"c9c002a8",
  1470 => x"a6e0c087",
  1471 => x"c078c048",
  1472 => x"e0c087c6",
  1473 => x"78c148a6",
  1474 => x"1e66e0c0",
  1475 => x"741ee0c0",
  1476 => x"c5d6ff49",
  1477 => x"d886c887",
  1478 => x"b7c058a6",
  1479 => x"dac106a8",
  1480 => x"8466d487",
  1481 => x"49bf66c4",
  1482 => x"7481e0c0",
  1483 => x"c3c14b89",
  1484 => x"fe714ac2",
  1485 => x"c287f9e5",
  1486 => x"4866dc84",
  1487 => x"e0c080c1",
  1488 => x"e4c058a6",
  1489 => x"81c14966",
  1490 => x"c002a970",
  1491 => x"e0c087c9",
  1492 => x"78c048a6",
  1493 => x"c087c6c0",
  1494 => x"c148a6e0",
  1495 => x"66e0c078",
  1496 => x"bf66c81e",
  1497 => x"81e0c049",
  1498 => x"1e718974",
  1499 => x"d4ff4974",
  1500 => x"86c887e8",
  1501 => x"01a8b7c0",
  1502 => x"dc87fefe",
  1503 => x"d0c00266",
  1504 => x"c9496e87",
  1505 => x"5166dc81",
  1506 => x"ccc1486e",
  1507 => x"ccc078f4",
  1508 => x"c9496e87",
  1509 => x"6e51c281",
  1510 => x"dad0c148",
  1511 => x"b766d078",
  1512 => x"c5c004ad",
  1513 => x"c085c187",
  1514 => x"66d087dc",
  1515 => x"d488c148",
  1516 => x"d1c058a6",
  1517 => x"cad3ff87",
  1518 => x"58a6d887",
  1519 => x"ff87c7c0",
  1520 => x"d887c0d3",
  1521 => x"66d458a6",
  1522 => x"87c9c002",
  1523 => x"b766c0c1",
  1524 => x"e4f504ad",
  1525 => x"adb7c787",
  1526 => x"87d9c003",
  1527 => x"91cb4975",
  1528 => x"8166f8c0",
  1529 => x"6a4aa1c4",
  1530 => x"7952c04a",
  1531 => x"b7c785c1",
  1532 => x"e7ff04ad",
  1533 => x"0266d887",
  1534 => x"c087e2c0",
  1535 => x"c14966f8",
  1536 => x"f8c081cd",
  1537 => x"d5c14a66",
  1538 => x"c152c082",
  1539 => x"c079d3cc",
  1540 => x"c14966f8",
  1541 => x"c3c181d1",
  1542 => x"d6c079c5",
  1543 => x"66f8c087",
  1544 => x"81cdc149",
  1545 => x"4a66f8c0",
  1546 => x"c182d1c1",
  1547 => x"c27accc3",
  1548 => x"c179f2c8",
  1549 => x"c04aebd0",
  1550 => x"c14966f8",
  1551 => x"797281d8",
  1552 => x"48bfd0ff",
  1553 => x"98c0c0c8",
  1554 => x"7058a6c4",
  1555 => x"d1c00298",
  1556 => x"bfd0ff87",
  1557 => x"c0c0c848",
  1558 => x"58a6c498",
  1559 => x"ff059870",
  1560 => x"d0ff87ef",
  1561 => x"78e0c048",
  1562 => x"ff4866cc",
  1563 => x"d2ff8ed8",
  1564 => x"c71e87da",
  1565 => x"c11ec01e",
  1566 => x"c21ef8e3",
  1567 => x"49bfece0",
  1568 => x"c187edef",
  1569 => x"c049f8e3",
  1570 => x"f487d4e6",
  1571 => x"1e4f268e",
  1572 => x"c287fdc9",
  1573 => x"c048c8e1",
  1574 => x"48d4ff50",
  1575 => x"c178ffc3",
  1576 => x"fe49d3c3",
  1577 => x"fe87e5df",
  1578 => x"7087f0e8",
  1579 => x"87cd0298",
  1580 => x"87edf4fe",
  1581 => x"c4029870",
  1582 => x"c24ac187",
  1583 => x"724ac087",
  1584 => x"87c8029a",
  1585 => x"49ddc3c1",
  1586 => x"87c0dffe",
  1587 => x"bff4e3c1",
  1588 => x"cbd6ff49",
  1589 => x"c0e1c287",
  1590 => x"c278c048",
  1591 => x"c048ece0",
  1592 => x"cdfe4978",
  1593 => x"87d4c387",
  1594 => x"c087f9c8",
  1595 => x"ff87d2e5",
  1596 => x"4f2687f6",
  1597 => x"000010e0",
  1598 => x"00001042",
  1599 => x"00002858",
  1600 => x"42000000",
  1601 => x"76000010",
  1602 => x"00000028",
  1603 => x"10420000",
  1604 => x"28940000",
  1605 => x"00000000",
  1606 => x"00104200",
  1607 => x"0028b200",
  1608 => x"00000000",
  1609 => x"00001042",
  1610 => x"000028d0",
  1611 => x"42000000",
  1612 => x"ee000010",
  1613 => x"00000028",
  1614 => x"10420000",
  1615 => x"290c0000",
  1616 => x"00000000",
  1617 => x"00131300",
  1618 => x"00000000",
  1619 => x"00000000",
  1620 => x"00001112",
  1621 => x"00000000",
  1622 => x"1e000000",
  1623 => x"87d5c11e",
  1624 => x"2658a6c4",
  1625 => x"711e4f26",
  1626 => x"48f0fe4a",
  1627 => x"0acd78c0",
  1628 => x"e5c10a7a",
  1629 => x"dcfe49fc",
  1630 => x"4f2687d2",
  1631 => x"20746553",
  1632 => x"646e6168",
  1633 => x"0a72656c",
  1634 => x"206e4900",
  1635 => x"65746e69",
  1636 => x"70757272",
  1637 => x"6f632074",
  1638 => x"7274736e",
  1639 => x"6f746375",
  1640 => x"1e000a72",
  1641 => x"49c9e6c1",
  1642 => x"87e0dbfe",
  1643 => x"49dbe5c1",
  1644 => x"2687f3fe",
  1645 => x"f0fe1e4f",
  1646 => x"4f2648bf",
  1647 => x"48f0fe1e",
  1648 => x"4f2678c1",
  1649 => x"48f0fe1e",
  1650 => x"4f2678c0",
  1651 => x"c04a711e",
  1652 => x"49a2c47a",
  1653 => x"a2c879c0",
  1654 => x"cc79c049",
  1655 => x"79c049a2",
  1656 => x"5e0e4f26",
  1657 => x"f80e5c5b",
  1658 => x"c84c7186",
  1659 => x"a4cc49a4",
  1660 => x"c1486b4b",
  1661 => x"58a6c480",
  1662 => x"a6c898cf",
  1663 => x"c4486958",
  1664 => x"d405a866",
  1665 => x"c1486b87",
  1666 => x"58a6c480",
  1667 => x"a6c898cf",
  1668 => x"c4486958",
  1669 => x"ec02a866",
  1670 => x"87e8fe87",
  1671 => x"49a4d0c1",
  1672 => x"90c4486b",
  1673 => x"7058a6c4",
  1674 => x"7966d481",
  1675 => x"80c1486b",
  1676 => x"cf58a6c8",
  1677 => x"c17b7098",
  1678 => x"fffd87d2",
  1679 => x"c28ef887",
  1680 => x"264d2687",
  1681 => x"264b264c",
  1682 => x"5b5e0e4f",
  1683 => x"f80e5d5c",
  1684 => x"c44d7186",
  1685 => x"486d4ca5",
  1686 => x"c505a86c",
  1687 => x"c048ff87",
  1688 => x"dffd87e5",
  1689 => x"4ba5d087",
  1690 => x"90c4486c",
  1691 => x"7058a6c4",
  1692 => x"c34b6b83",
  1693 => x"486c9bff",
  1694 => x"a6c880c1",
  1695 => x"7098cf58",
  1696 => x"87f8fc7c",
  1697 => x"f8484973",
  1698 => x"87f5fe8e",
  1699 => x"f81e731e",
  1700 => x"87f0fc86",
  1701 => x"494bbfe0",
  1702 => x"99c0e0c0",
  1703 => x"87e7c002",
  1704 => x"ffc34a73",
  1705 => x"eae4c29a",
  1706 => x"90c448bf",
  1707 => x"c258a6c4",
  1708 => x"7049fae4",
  1709 => x"c2797281",
  1710 => x"48bfeae4",
  1711 => x"a6c880c1",
  1712 => x"c298cf58",
  1713 => x"7358eee4",
  1714 => x"99c0d049",
  1715 => x"87f2c002",
  1716 => x"bff2e4c2",
  1717 => x"f6e4c248",
  1718 => x"c002a8bf",
  1719 => x"e4c287e4",
  1720 => x"c448bff2",
  1721 => x"58a6c490",
  1722 => x"49fae5c2",
  1723 => x"48e08170",
  1724 => x"e4c27869",
  1725 => x"c148bff2",
  1726 => x"58a6c880",
  1727 => x"e4c298cf",
  1728 => x"f0fa58f6",
  1729 => x"58a6c487",
  1730 => x"f887f1fa",
  1731 => x"87f5fc8e",
  1732 => x"eae4c21e",
  1733 => x"87f4fa49",
  1734 => x"49cceac1",
  1735 => x"c387c7f9",
  1736 => x"4f2687f5",
  1737 => x"c21e731e",
  1738 => x"fc49eae4",
  1739 => x"4a7087db",
  1740 => x"04aab7c0",
  1741 => x"c387ccc2",
  1742 => x"c905aaf0",
  1743 => x"cfefc187",
  1744 => x"c178c148",
  1745 => x"e0c387ed",
  1746 => x"87c905aa",
  1747 => x"48d3efc1",
  1748 => x"dec178c1",
  1749 => x"d3efc187",
  1750 => x"87c602bf",
  1751 => x"4ba2c0c2",
  1752 => x"4b7287c2",
  1753 => x"bfcfefc1",
  1754 => x"87e0c002",
  1755 => x"b7c44973",
  1756 => x"efc19129",
  1757 => x"4a7381d7",
  1758 => x"92c29acf",
  1759 => x"307248c1",
  1760 => x"baff4a70",
  1761 => x"98694872",
  1762 => x"87db7970",
  1763 => x"b7c44973",
  1764 => x"efc19129",
  1765 => x"4a7381d7",
  1766 => x"92c29acf",
  1767 => x"307248c3",
  1768 => x"69484a70",
  1769 => x"c17970b0",
  1770 => x"c048d3ef",
  1771 => x"cfefc178",
  1772 => x"c278c048",
  1773 => x"fa49eae4",
  1774 => x"4a7087cf",
  1775 => x"03aab7c0",
  1776 => x"c087f4fd",
  1777 => x"2687c448",
  1778 => x"264c264d",
  1779 => x"004f264b",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"1e000000",
  1798 => x"49724ac0",
  1799 => x"efc191c4",
  1800 => x"79c081d7",
  1801 => x"b7d082c1",
  1802 => x"87ee04aa",
  1803 => x"5e0e4f26",
  1804 => x"0e5d5c5b",
  1805 => x"cbf64d71",
  1806 => x"c44a7587",
  1807 => x"c1922ab7",
  1808 => x"7582d7ef",
  1809 => x"c29ccf4c",
  1810 => x"4b496a94",
  1811 => x"9bc32b74",
  1812 => x"307448c2",
  1813 => x"bcff4c70",
  1814 => x"98714874",
  1815 => x"dbf57a70",
  1816 => x"fd487387",
  1817 => x"1e1e87e1",
  1818 => x"48bfd0ff",
  1819 => x"98c0c0c8",
  1820 => x"7058a6c4",
  1821 => x"87d00298",
  1822 => x"48bfd0ff",
  1823 => x"98c0c0c8",
  1824 => x"7058a6c4",
  1825 => x"87f00598",
  1826 => x"c448d0ff",
  1827 => x"487178e1",
  1828 => x"7808d4ff",
  1829 => x"ff4866c8",
  1830 => x"267808d4",
  1831 => x"1e1e4f26",
  1832 => x"66c84a71",
  1833 => x"49721e49",
  1834 => x"c487fbfe",
  1835 => x"bfd0ff86",
  1836 => x"c0c0c848",
  1837 => x"58a6c498",
  1838 => x"d0029870",
  1839 => x"bfd0ff87",
  1840 => x"c0c0c848",
  1841 => x"58a6c498",
  1842 => x"f0059870",
  1843 => x"48d0ff87",
  1844 => x"2678e0c0",
  1845 => x"731e4f26",
  1846 => x"c84b711e",
  1847 => x"4a731e66",
  1848 => x"49a2e0c1",
  1849 => x"2687f7fe",
  1850 => x"4d2687c4",
  1851 => x"4b264c26",
  1852 => x"1e1e4f26",
  1853 => x"48bfd0ff",
  1854 => x"98c0c0c8",
  1855 => x"7058a6c4",
  1856 => x"87d00298",
  1857 => x"48bfd0ff",
  1858 => x"98c0c0c8",
  1859 => x"7058a6c4",
  1860 => x"87f00598",
  1861 => x"c448d0ff",
  1862 => x"487178c9",
  1863 => x"7808d4ff",
  1864 => x"1e4f2626",
  1865 => x"494a711e",
  1866 => x"ff87c7ff",
  1867 => x"c848bfd0",
  1868 => x"c498c0c0",
  1869 => x"987058a6",
  1870 => x"ff87d002",
  1871 => x"c848bfd0",
  1872 => x"c498c0c0",
  1873 => x"987058a6",
  1874 => x"ff87f005",
  1875 => x"78c848d0",
  1876 => x"1e4f2626",
  1877 => x"711e1e73",
  1878 => x"c6e7c24b",
  1879 => x"87c302bf",
  1880 => x"ff87ccc3",
  1881 => x"c848bfd0",
  1882 => x"c498c0c0",
  1883 => x"987058a6",
  1884 => x"ff87d002",
  1885 => x"c848bfd0",
  1886 => x"c498c0c0",
  1887 => x"987058a6",
  1888 => x"ff87f005",
  1889 => x"c9c448d0",
  1890 => x"c0487378",
  1891 => x"d4ffb0e0",
  1892 => x"e6c27808",
  1893 => x"78c048fa",
  1894 => x"c50266cc",
  1895 => x"49ffc387",
  1896 => x"49c087c2",
  1897 => x"59c2e7c2",
  1898 => x"c60266d0",
  1899 => x"d5d5c587",
  1900 => x"cf87c44a",
  1901 => x"c24affff",
  1902 => x"c25ac6e7",
  1903 => x"c148c6e7",
  1904 => x"87c42678",
  1905 => x"4c264d26",
  1906 => x"4f264b26",
  1907 => x"5c5b5e0e",
  1908 => x"4a710e5d",
  1909 => x"bfc2e7c2",
  1910 => x"029a724c",
  1911 => x"c84987cb",
  1912 => x"cdf6c191",
  1913 => x"c483714b",
  1914 => x"cdfac187",
  1915 => x"134dc04b",
  1916 => x"c2997449",
  1917 => x"48bffee6",
  1918 => x"d4ffb871",
  1919 => x"b7c17808",
  1920 => x"b7c8852c",
  1921 => x"87e704ad",
  1922 => x"bffae6c2",
  1923 => x"c280c848",
  1924 => x"fe58fee6",
  1925 => x"731e87ee",
  1926 => x"134b711e",
  1927 => x"cb029a4a",
  1928 => x"fe497287",
  1929 => x"4a1387e6",
  1930 => x"87f5059a",
  1931 => x"1e87d9fe",
  1932 => x"fae6c21e",
  1933 => x"e6c249bf",
  1934 => x"a1c148fa",
  1935 => x"b7c0c478",
  1936 => x"87db03a9",
  1937 => x"c248d4ff",
  1938 => x"78bffee6",
  1939 => x"bffae6c2",
  1940 => x"fae6c249",
  1941 => x"78a1c148",
  1942 => x"a9b7c0c4",
  1943 => x"ff87e504",
  1944 => x"c848bfd0",
  1945 => x"c498c0c0",
  1946 => x"987058a6",
  1947 => x"ff87d002",
  1948 => x"c848bfd0",
  1949 => x"c498c0c0",
  1950 => x"987058a6",
  1951 => x"ff87f005",
  1952 => x"78c848d0",
  1953 => x"48c6e7c2",
  1954 => x"262678c0",
  1955 => x"0000004f",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00005f5f",
  1959 => x"03030000",
  1960 => x"00030300",
  1961 => x"7f7f1400",
  1962 => x"147f7f14",
  1963 => x"2e240000",
  1964 => x"123a6b6b",
  1965 => x"366a4c00",
  1966 => x"32566c18",
  1967 => x"4f7e3000",
  1968 => x"683a7759",
  1969 => x"04000040",
  1970 => x"00000307",
  1971 => x"1c000000",
  1972 => x"0041633e",
  1973 => x"41000000",
  1974 => x"001c3e63",
  1975 => x"3e2a0800",
  1976 => x"2a3e1c1c",
  1977 => x"08080008",
  1978 => x"08083e3e",
  1979 => x"80000000",
  1980 => x"000060e0",
  1981 => x"08080000",
  1982 => x"08080808",
  1983 => x"00000000",
  1984 => x"00006060",
  1985 => x"30604000",
  1986 => x"03060c18",
  1987 => x"7f3e0001",
  1988 => x"3e7f4d59",
  1989 => x"06040000",
  1990 => x"00007f7f",
  1991 => x"63420000",
  1992 => x"464f5971",
  1993 => x"63220000",
  1994 => x"367f4949",
  1995 => x"161c1800",
  1996 => x"107f7f13",
  1997 => x"67270000",
  1998 => x"397d4545",
  1999 => x"7e3c0000",
  2000 => x"3079494b",
  2001 => x"01010000",
  2002 => x"070f7971",
  2003 => x"7f360000",
  2004 => x"367f4949",
  2005 => x"4f060000",
  2006 => x"1e3f6949",
  2007 => x"00000000",
  2008 => x"00006666",
  2009 => x"80000000",
  2010 => x"000066e6",
  2011 => x"08080000",
  2012 => x"22221414",
  2013 => x"14140000",
  2014 => x"14141414",
  2015 => x"22220000",
  2016 => x"08081414",
  2017 => x"03020000",
  2018 => x"060f5951",
  2019 => x"417f3e00",
  2020 => x"1e1f555d",
  2021 => x"7f7e0000",
  2022 => x"7e7f0909",
  2023 => x"7f7f0000",
  2024 => x"367f4949",
  2025 => x"3e1c0000",
  2026 => x"41414163",
  2027 => x"7f7f0000",
  2028 => x"1c3e6341",
  2029 => x"7f7f0000",
  2030 => x"41414949",
  2031 => x"7f7f0000",
  2032 => x"01010909",
  2033 => x"7f3e0000",
  2034 => x"7a7b4941",
  2035 => x"7f7f0000",
  2036 => x"7f7f0808",
  2037 => x"41000000",
  2038 => x"00417f7f",
  2039 => x"60200000",
  2040 => x"3f7f4040",
  2041 => x"087f7f00",
  2042 => x"4163361c",
  2043 => x"7f7f0000",
  2044 => x"40404040",
  2045 => x"067f7f00",
  2046 => x"7f7f060c",
  2047 => x"067f7f00",
  2048 => x"7f7f180c",
  2049 => x"7f3e0000",
  2050 => x"3e7f4141",
  2051 => x"7f7f0000",
  2052 => x"060f0909",
  2053 => x"417f3e00",
  2054 => x"407e7f61",
  2055 => x"7f7f0000",
  2056 => x"667f1909",
  2057 => x"6f260000",
  2058 => x"327b594d",
  2059 => x"01010000",
  2060 => x"01017f7f",
  2061 => x"7f3f0000",
  2062 => x"3f7f4040",
  2063 => x"3f0f0000",
  2064 => x"0f3f7070",
  2065 => x"307f7f00",
  2066 => x"7f7f3018",
  2067 => x"36634100",
  2068 => x"63361c1c",
  2069 => x"06030141",
  2070 => x"03067c7c",
  2071 => x"59716101",
  2072 => x"4143474d",
  2073 => x"7f000000",
  2074 => x"0041417f",
  2075 => x"06030100",
  2076 => x"6030180c",
  2077 => x"41000040",
  2078 => x"007f7f41",
  2079 => x"060c0800",
  2080 => x"080c0603",
  2081 => x"80808000",
  2082 => x"80808080",
  2083 => x"00000000",
  2084 => x"00040703",
  2085 => x"74200000",
  2086 => x"787c5454",
  2087 => x"7f7f0000",
  2088 => x"387c4444",
  2089 => x"7c380000",
  2090 => x"00444444",
  2091 => x"7c380000",
  2092 => x"7f7f4444",
  2093 => x"7c380000",
  2094 => x"185c5454",
  2095 => x"7e040000",
  2096 => x"0005057f",
  2097 => x"bc180000",
  2098 => x"7cfca4a4",
  2099 => x"7f7f0000",
  2100 => x"787c0404",
  2101 => x"00000000",
  2102 => x"00407d3d",
  2103 => x"80800000",
  2104 => x"007dfd80",
  2105 => x"7f7f0000",
  2106 => x"446c3810",
  2107 => x"00000000",
  2108 => x"00407f3f",
  2109 => x"0c7c7c00",
  2110 => x"787c0c18",
  2111 => x"7c7c0000",
  2112 => x"787c0404",
  2113 => x"7c380000",
  2114 => x"387c4444",
  2115 => x"fcfc0000",
  2116 => x"183c2424",
  2117 => x"3c180000",
  2118 => x"fcfc2424",
  2119 => x"7c7c0000",
  2120 => x"080c0404",
  2121 => x"5c480000",
  2122 => x"20745454",
  2123 => x"3f040000",
  2124 => x"0044447f",
  2125 => x"7c3c0000",
  2126 => x"7c7c4040",
  2127 => x"3c1c0000",
  2128 => x"1c3c6060",
  2129 => x"607c3c00",
  2130 => x"3c7c6030",
  2131 => x"386c4400",
  2132 => x"446c3810",
  2133 => x"bc1c0000",
  2134 => x"1c3c60e0",
  2135 => x"64440000",
  2136 => x"444c5c74",
  2137 => x"08080000",
  2138 => x"4141773e",
  2139 => x"00000000",
  2140 => x"00007f7f",
  2141 => x"41410000",
  2142 => x"08083e77",
  2143 => x"01010200",
  2144 => x"01020203",
  2145 => x"7f7f7f00",
  2146 => x"7f7f7f7f",
  2147 => x"1c080800",
  2148 => x"7f3e3e1c",
  2149 => x"3e7f7f7f",
  2150 => x"081c1c3e",
  2151 => x"18100008",
  2152 => x"10187c7c",
  2153 => x"30100000",
  2154 => x"10307c7c",
  2155 => x"60301000",
  2156 => x"061e7860",
  2157 => x"3c664200",
  2158 => x"42663c18",
  2159 => x"6a387800",
  2160 => x"386cc6c2",
  2161 => x"00006000",
  2162 => x"60000060",
  2163 => x"5b5e0e00",
  2164 => x"1e0e5d5c",
  2165 => x"e7c24c71",
  2166 => x"c04dbfce",
  2167 => x"741ec04b",
  2168 => x"87c702ab",
  2169 => x"c048a6c4",
  2170 => x"c487c578",
  2171 => x"78c148a6",
  2172 => x"731e66c4",
  2173 => x"87dbed49",
  2174 => x"e0c086c8",
  2175 => x"87ccef49",
  2176 => x"6a4aa5c4",
  2177 => x"87cef049",
  2178 => x"cb87e4f0",
  2179 => x"c883c185",
  2180 => x"ff04abb7",
  2181 => x"262687c7",
  2182 => x"264c264d",
  2183 => x"1e4f264b",
  2184 => x"e7c24a71",
  2185 => x"e7c25ad2",
  2186 => x"78c748d2",
  2187 => x"87ddfe49",
  2188 => x"c11e4f26",
  2189 => x"eaeb49c0",
  2190 => x"e2d2c287",
  2191 => x"2678c048",
  2192 => x"5b5e0e4f",
  2193 => x"f40e5d5c",
  2194 => x"c87ec086",
  2195 => x"bfec48a6",
  2196 => x"c280fc78",
  2197 => x"78bfcee7",
  2198 => x"bfd6e7c2",
  2199 => x"4cbfe84d",
  2200 => x"c9e749c7",
  2201 => x"c2497087",
  2202 => x"87d00599",
  2203 => x"bfdad2c2",
  2204 => x"c8b9ff49",
  2205 => x"99c19966",
  2206 => x"87ebc002",
  2207 => x"ede649c7",
  2208 => x"02987087",
  2209 => x"dbe287cd",
  2210 => x"e649c787",
  2211 => x"987087e0",
  2212 => x"c287f305",
  2213 => x"4abfe2d2",
  2214 => x"d2c2bac1",
  2215 => x"c0c15ae6",
  2216 => x"fee949a2",
  2217 => x"c27ec187",
  2218 => x"c848dad2",
  2219 => x"d2c27866",
  2220 => x"c105bfe2",
  2221 => x"c0c887cb",
  2222 => x"d2c27ec0",
  2223 => x"49134bca",
  2224 => x"7087ebe5",
  2225 => x"87c20298",
  2226 => x"486eb46e",
  2227 => x"c428b7c1",
  2228 => x"987058a6",
  2229 => x"87e6ff05",
  2230 => x"ffc34974",
  2231 => x"c01e7199",
  2232 => x"87f2e749",
  2233 => x"b7c84974",
  2234 => x"c11e7129",
  2235 => x"87e6e749",
  2236 => x"fdc386c8",
  2237 => x"87f6e449",
  2238 => x"e449fac3",
  2239 => x"c4c687f0",
  2240 => x"c3497487",
  2241 => x"b7c899ff",
  2242 => x"74b4712c",
  2243 => x"e2c0029c",
  2244 => x"48a6c887",
  2245 => x"78bfc8ff",
  2246 => x"c24966c8",
  2247 => x"89bfded2",
  2248 => x"03a9c0c2",
  2249 => x"4cc087c4",
  2250 => x"d2c287cf",
  2251 => x"66c848de",
  2252 => x"c287c678",
  2253 => x"c048ded2",
  2254 => x"c8497478",
  2255 => x"87ce0599",
  2256 => x"e349f5c3",
  2257 => x"497087e8",
  2258 => x"c00299c2",
  2259 => x"e7c287e6",
  2260 => x"c902bfd2",
  2261 => x"88c14887",
  2262 => x"58d6e7c2",
  2263 => x"66c487d4",
  2264 => x"80d8c148",
  2265 => x"6e58a6c4",
  2266 => x"c5c002bf",
  2267 => x"49ff4b87",
  2268 => x"7ec10f73",
  2269 => x"99c44974",
  2270 => x"c387ce05",
  2271 => x"ede249f2",
  2272 => x"c2497087",
  2273 => x"eec00299",
  2274 => x"d2e7c287",
  2275 => x"486e7ebf",
  2276 => x"03a8b7c7",
  2277 => x"6e87cac0",
  2278 => x"c280c148",
  2279 => x"d458d6e7",
  2280 => x"4866c487",
  2281 => x"c480d8c1",
  2282 => x"bf6e58a6",
  2283 => x"87c5c002",
  2284 => x"7349fe4b",
  2285 => x"c37ec10f",
  2286 => x"f1e149fd",
  2287 => x"c2497087",
  2288 => x"e3c00299",
  2289 => x"d2e7c287",
  2290 => x"c9c002bf",
  2291 => x"d2e7c287",
  2292 => x"c078c048",
  2293 => x"66c487d0",
  2294 => x"82d8c14a",
  2295 => x"c5c0026a",
  2296 => x"49fd4b87",
  2297 => x"7ec10f73",
  2298 => x"e149fac3",
  2299 => x"497087c0",
  2300 => x"c00299c2",
  2301 => x"e7c287eb",
  2302 => x"c748bfd2",
  2303 => x"c003a8b7",
  2304 => x"e7c287c9",
  2305 => x"78c748d2",
  2306 => x"c487d4c0",
  2307 => x"d8c14866",
  2308 => x"58a6c480",
  2309 => x"c002bf6e",
  2310 => x"fc4b87c5",
  2311 => x"c10f7349",
  2312 => x"c349747e",
  2313 => x"c00599f0",
  2314 => x"dac187cf",
  2315 => x"fddfff49",
  2316 => x"c2497087",
  2317 => x"d0c00299",
  2318 => x"d2e7c287",
  2319 => x"cb4b49bf",
  2320 => x"8366c493",
  2321 => x"73714b6b",
  2322 => x"029d750f",
  2323 => x"6d87e9c0",
  2324 => x"87e4c002",
  2325 => x"dfff496d",
  2326 => x"497087d4",
  2327 => x"c00299c1",
  2328 => x"a5c487cb",
  2329 => x"d2e7c24b",
  2330 => x"4b6b49bf",
  2331 => x"0285c80f",
  2332 => x"6d87c5c0",
  2333 => x"87dcff05",
  2334 => x"c8c0026e",
  2335 => x"d2e7c287",
  2336 => x"c8f549bf",
  2337 => x"f68ef487",
  2338 => x"125887cd",
  2339 => x"1b1d1411",
  2340 => x"595a231c",
  2341 => x"f2f59491",
  2342 => x"0000f4eb",
  2343 => x"00000000",
  2344 => x"00000000",
  2345 => x"19a30000",
  2346 => x"19a30000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
