
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"c4",x"c3",x"87"),
    12 => (x"86",x"c0",x"d0",x"4e"),
    13 => (x"49",x"f4",x"c4",x"c3"),
    14 => (x"48",x"c4",x"f0",x"c2"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"c4",x"f0",x"c2",x"87"),
    21 => (x"c0",x"f0",x"c2",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"f7",x"c1",x"87",x"f7"),
    25 => (x"f0",x"c2",x"87",x"fe"),
    26 => (x"f0",x"c2",x"4d",x"c4"),
    27 => (x"ad",x"74",x"4c",x"c4"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"5c",x"5b",x"5e",x"0e"),
    32 => (x"86",x"f0",x"0e",x"5d"),
    33 => (x"a6",x"c4",x"4c",x"c0"),
    34 => (x"c0",x"78",x"c0",x"48"),
    35 => (x"c0",x"4b",x"a6",x"e4"),
    36 => (x"48",x"49",x"66",x"e0"),
    37 => (x"e4",x"c0",x"80",x"c1"),
    38 => (x"48",x"11",x"58",x"a6"),
    39 => (x"70",x"58",x"a6",x"c4"),
    40 => (x"f6",x"c3",x"02",x"98"),
    41 => (x"02",x"66",x"c4",x"87"),
    42 => (x"c4",x"87",x"c6",x"c3"),
    43 => (x"78",x"c0",x"48",x"a6"),
    44 => (x"f0",x"c0",x"4a",x"6e"),
    45 => (x"da",x"c2",x"02",x"8a"),
    46 => (x"8a",x"f3",x"c0",x"87"),
    47 => (x"87",x"db",x"c2",x"02"),
    48 => (x"dc",x"02",x"8a",x"c1"),
    49 => (x"02",x"8a",x"c8",x"87"),
    50 => (x"c4",x"87",x"c8",x"c2"),
    51 => (x"87",x"d1",x"02",x"8a"),
    52 => (x"c1",x"02",x"8a",x"c3"),
    53 => (x"8a",x"c2",x"87",x"eb"),
    54 => (x"c3",x"87",x"c6",x"02"),
    55 => (x"c9",x"c2",x"05",x"8a"),
    56 => (x"73",x"83",x"c4",x"87"),
    57 => (x"69",x"89",x"c4",x"49"),
    58 => (x"c1",x"02",x"6e",x"7e"),
    59 => (x"a6",x"c8",x"87",x"c8"),
    60 => (x"c4",x"78",x"c0",x"48"),
    61 => (x"cc",x"78",x"c0",x"80"),
    62 => (x"4a",x"6e",x"4d",x"66"),
    63 => (x"cf",x"2a",x"b7",x"dc"),
    64 => (x"c4",x"48",x"6e",x"9a"),
    65 => (x"72",x"58",x"a6",x"30"),
    66 => (x"87",x"c5",x"02",x"9a"),
    67 => (x"c1",x"48",x"a6",x"c8"),
    68 => (x"06",x"aa",x"c9",x"78"),
    69 => (x"f7",x"c0",x"87",x"c5"),
    70 => (x"c0",x"87",x"c3",x"82"),
    71 => (x"66",x"c8",x"82",x"f0"),
    72 => (x"72",x"87",x"c7",x"02"),
    73 => (x"87",x"f3",x"c2",x"49"),
    74 => (x"85",x"c1",x"84",x"c1"),
    75 => (x"04",x"ad",x"b7",x"c8"),
    76 => (x"c1",x"87",x"c7",x"ff"),
    77 => (x"f0",x"c0",x"87",x"cf"),
    78 => (x"87",x"df",x"c2",x"49"),
    79 => (x"c4",x"c1",x"84",x"c1"),
    80 => (x"73",x"83",x"c4",x"87"),
    81 => (x"6a",x"8a",x"c4",x"4a"),
    82 => (x"87",x"db",x"c1",x"49"),
    83 => (x"4c",x"a4",x"49",x"70"),
    84 => (x"c4",x"87",x"f2",x"c0"),
    85 => (x"78",x"c1",x"48",x"a6"),
    86 => (x"c4",x"87",x"ea",x"c0"),
    87 => (x"c4",x"4a",x"73",x"83"),
    88 => (x"c1",x"49",x"6a",x"8a"),
    89 => (x"84",x"c1",x"87",x"f5"),
    90 => (x"49",x"6e",x"87",x"db"),
    91 => (x"d4",x"87",x"ec",x"c1"),
    92 => (x"c0",x"48",x"6e",x"87"),
    93 => (x"c7",x"05",x"a8",x"e5"),
    94 => (x"48",x"a6",x"c4",x"87"),
    95 => (x"87",x"c5",x"78",x"c1"),
    96 => (x"d6",x"c1",x"49",x"6e"),
    97 => (x"66",x"e0",x"c0",x"87"),
    98 => (x"80",x"c1",x"48",x"49"),
    99 => (x"58",x"a6",x"e4",x"c0"),
   100 => (x"a6",x"c4",x"48",x"11"),
   101 => (x"05",x"98",x"70",x"58"),
   102 => (x"74",x"87",x"ca",x"fc"),
   103 => (x"26",x"8e",x"f0",x"48"),
   104 => (x"26",x"4c",x"26",x"4d"),
   105 => (x"0e",x"4f",x"26",x"4b"),
   106 => (x"0e",x"5c",x"5b",x"5e"),
   107 => (x"4c",x"c0",x"4b",x"71"),
   108 => (x"02",x"9a",x"4a",x"13"),
   109 => (x"49",x"72",x"87",x"cd"),
   110 => (x"c1",x"87",x"e0",x"c0"),
   111 => (x"9a",x"4a",x"13",x"84"),
   112 => (x"74",x"87",x"f3",x"05"),
   113 => (x"26",x"4c",x"26",x"48"),
   114 => (x"1e",x"4f",x"26",x"4b"),
   115 => (x"73",x"81",x"48",x"73"),
   116 => (x"87",x"c5",x"02",x"a9"),
   117 => (x"f6",x"05",x"53",x"12"),
   118 => (x"1e",x"4f",x"26",x"87"),
   119 => (x"4a",x"c0",x"ff",x"1e"),
   120 => (x"c0",x"c4",x"48",x"6a"),
   121 => (x"58",x"a6",x"c4",x"98"),
   122 => (x"f3",x"02",x"98",x"70"),
   123 => (x"48",x"7a",x"71",x"87"),
   124 => (x"1e",x"4f",x"26",x"26"),
   125 => (x"d4",x"ff",x"1e",x"73"),
   126 => (x"7b",x"ff",x"c3",x"4b"),
   127 => (x"ff",x"c3",x"4a",x"6b"),
   128 => (x"c8",x"49",x"6b",x"7b"),
   129 => (x"c3",x"b1",x"72",x"32"),
   130 => (x"4a",x"6b",x"7b",x"ff"),
   131 => (x"b2",x"71",x"31",x"c8"),
   132 => (x"6b",x"7b",x"ff",x"c3"),
   133 => (x"72",x"32",x"c8",x"49"),
   134 => (x"c4",x"48",x"71",x"b1"),
   135 => (x"26",x"4d",x"26",x"87"),
   136 => (x"26",x"4b",x"26",x"4c"),
   137 => (x"5b",x"5e",x"0e",x"4f"),
   138 => (x"71",x"0e",x"5d",x"5c"),
   139 => (x"4c",x"d4",x"ff",x"4a"),
   140 => (x"ff",x"c3",x"48",x"72"),
   141 => (x"c2",x"7c",x"70",x"98"),
   142 => (x"05",x"bf",x"c4",x"f0"),
   143 => (x"66",x"d0",x"87",x"c8"),
   144 => (x"d4",x"30",x"c9",x"48"),
   145 => (x"66",x"d0",x"58",x"a6"),
   146 => (x"71",x"29",x"d8",x"49"),
   147 => (x"98",x"ff",x"c3",x"48"),
   148 => (x"66",x"d0",x"7c",x"70"),
   149 => (x"71",x"29",x"d0",x"49"),
   150 => (x"98",x"ff",x"c3",x"48"),
   151 => (x"66",x"d0",x"7c",x"70"),
   152 => (x"71",x"29",x"c8",x"49"),
   153 => (x"98",x"ff",x"c3",x"48"),
   154 => (x"66",x"d0",x"7c",x"70"),
   155 => (x"98",x"ff",x"c3",x"48"),
   156 => (x"49",x"72",x"7c",x"70"),
   157 => (x"48",x"71",x"29",x"d0"),
   158 => (x"70",x"98",x"ff",x"c3"),
   159 => (x"c9",x"4b",x"6c",x"7c"),
   160 => (x"c3",x"4d",x"ff",x"f0"),
   161 => (x"d0",x"05",x"ab",x"ff"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"8d",x"c1",x"4b",x"6c"),
   164 => (x"c3",x"87",x"c6",x"02"),
   165 => (x"f0",x"02",x"ab",x"ff"),
   166 => (x"fd",x"48",x"73",x"87"),
   167 => (x"c0",x"1e",x"87",x"ff"),
   168 => (x"48",x"d4",x"ff",x"49"),
   169 => (x"c1",x"78",x"ff",x"c3"),
   170 => (x"b7",x"c8",x"c3",x"81"),
   171 => (x"87",x"f1",x"04",x"a9"),
   172 => (x"73",x"1e",x"4f",x"26"),
   173 => (x"c4",x"87",x"e7",x"1e"),
   174 => (x"c0",x"4b",x"df",x"f8"),
   175 => (x"f0",x"ff",x"c0",x"1e"),
   176 => (x"fd",x"49",x"f7",x"c1"),
   177 => (x"86",x"c4",x"87",x"df"),
   178 => (x"c0",x"05",x"a8",x"c1"),
   179 => (x"d4",x"ff",x"87",x"ea"),
   180 => (x"78",x"ff",x"c3",x"48"),
   181 => (x"c0",x"c0",x"c0",x"c1"),
   182 => (x"c0",x"1e",x"c0",x"c0"),
   183 => (x"e9",x"c1",x"f0",x"e1"),
   184 => (x"87",x"c1",x"fd",x"49"),
   185 => (x"98",x"70",x"86",x"c4"),
   186 => (x"ff",x"87",x"ca",x"05"),
   187 => (x"ff",x"c3",x"48",x"d4"),
   188 => (x"cb",x"48",x"c1",x"78"),
   189 => (x"87",x"e6",x"fe",x"87"),
   190 => (x"fe",x"05",x"8b",x"c1"),
   191 => (x"48",x"c0",x"87",x"fd"),
   192 => (x"1e",x"87",x"de",x"fc"),
   193 => (x"d4",x"ff",x"1e",x"73"),
   194 => (x"78",x"ff",x"c3",x"48"),
   195 => (x"fa",x"49",x"fe",x"cc"),
   196 => (x"4b",x"d3",x"87",x"d5"),
   197 => (x"ff",x"c0",x"1e",x"c0"),
   198 => (x"49",x"c1",x"c1",x"f0"),
   199 => (x"c4",x"87",x"c6",x"fc"),
   200 => (x"05",x"98",x"70",x"86"),
   201 => (x"d4",x"ff",x"87",x"ca"),
   202 => (x"78",x"ff",x"c3",x"48"),
   203 => (x"87",x"cb",x"48",x"c1"),
   204 => (x"c1",x"87",x"eb",x"fd"),
   205 => (x"db",x"ff",x"05",x"8b"),
   206 => (x"fb",x"48",x"c0",x"87"),
   207 => (x"4d",x"43",x"87",x"e3"),
   208 => (x"4d",x"43",x"00",x"44"),
   209 => (x"20",x"38",x"35",x"44"),
   210 => (x"20",x"0a",x"64",x"25"),
   211 => (x"4d",x"43",x"00",x"20"),
   212 => (x"5f",x"38",x"35",x"44"),
   213 => (x"64",x"25",x"20",x"32"),
   214 => (x"00",x"20",x"20",x"0a"),
   215 => (x"35",x"44",x"4d",x"43"),
   216 => (x"64",x"25",x"20",x"38"),
   217 => (x"00",x"20",x"20",x"0a"),
   218 => (x"43",x"48",x"44",x"53"),
   219 => (x"69",x"6e",x"49",x"20"),
   220 => (x"6c",x"61",x"69",x"74"),
   221 => (x"74",x"61",x"7a",x"69"),
   222 => (x"20",x"6e",x"6f",x"69"),
   223 => (x"6f",x"72",x"72",x"65"),
   224 => (x"00",x"0a",x"21",x"72"),
   225 => (x"5f",x"64",x"6d",x"63"),
   226 => (x"38",x"44",x"4d",x"43"),
   227 => (x"73",x"65",x"72",x"20"),
   228 => (x"73",x"6e",x"6f",x"70"),
   229 => (x"25",x"20",x"3a",x"65"),
   230 => (x"49",x"00",x"0a",x"64"),
   231 => (x"00",x"52",x"52",x"45"),
   232 => (x"00",x"49",x"50",x"53"),
   233 => (x"63",x"20",x"44",x"53"),
   234 => (x"20",x"64",x"72",x"61"),
   235 => (x"65",x"7a",x"69",x"73"),
   236 => (x"20",x"73",x"69",x"20"),
   237 => (x"00",x"0a",x"64",x"25"),
   238 => (x"74",x"69",x"72",x"57"),
   239 => (x"61",x"66",x"20",x"65"),
   240 => (x"64",x"65",x"6c",x"69"),
   241 => (x"5f",x"63",x"00",x"0a"),
   242 => (x"65",x"7a",x"69",x"73"),
   243 => (x"6c",x"75",x"6d",x"5f"),
   244 => (x"25",x"20",x"3a",x"74"),
   245 => (x"72",x"20",x"2c",x"64"),
   246 => (x"5f",x"64",x"61",x"65"),
   247 => (x"6c",x"5f",x"6c",x"62"),
   248 => (x"20",x"3a",x"6e",x"65"),
   249 => (x"20",x"2c",x"64",x"25"),
   250 => (x"7a",x"69",x"73",x"63"),
   251 => (x"25",x"20",x"3a",x"65"),
   252 => (x"4d",x"00",x"0a",x"64"),
   253 => (x"20",x"74",x"6c",x"75"),
   254 => (x"00",x"0a",x"64",x"25"),
   255 => (x"62",x"20",x"64",x"25"),
   256 => (x"6b",x"63",x"6f",x"6c"),
   257 => (x"66",x"6f",x"20",x"73"),
   258 => (x"7a",x"69",x"73",x"20"),
   259 => (x"64",x"25",x"20",x"65"),
   260 => (x"64",x"25",x"00",x"0a"),
   261 => (x"6f",x"6c",x"62",x"20"),
   262 => (x"20",x"73",x"6b",x"63"),
   263 => (x"35",x"20",x"66",x"6f"),
   264 => (x"62",x"20",x"32",x"31"),
   265 => (x"73",x"65",x"74",x"79"),
   266 => (x"5e",x"0e",x"00",x"0a"),
   267 => (x"0e",x"5d",x"5c",x"5b"),
   268 => (x"f9",x"4d",x"d4",x"ff"),
   269 => (x"ea",x"c6",x"87",x"e8"),
   270 => (x"f0",x"e1",x"c0",x"1e"),
   271 => (x"f7",x"49",x"c8",x"c1"),
   272 => (x"4b",x"70",x"87",x"e3"),
   273 => (x"1e",x"c4",x"ce",x"1e"),
   274 => (x"cc",x"87",x"f1",x"f0"),
   275 => (x"02",x"ab",x"c1",x"86"),
   276 => (x"ee",x"fa",x"87",x"c8"),
   277 => (x"c2",x"48",x"c0",x"87"),
   278 => (x"d6",x"f6",x"87",x"ca"),
   279 => (x"cf",x"49",x"70",x"87"),
   280 => (x"c6",x"99",x"ff",x"ff"),
   281 => (x"c8",x"02",x"a9",x"ea"),
   282 => (x"87",x"d7",x"fa",x"87"),
   283 => (x"f3",x"c1",x"48",x"c0"),
   284 => (x"7d",x"ff",x"c3",x"87"),
   285 => (x"f8",x"4c",x"f1",x"c0"),
   286 => (x"98",x"70",x"87",x"f8"),
   287 => (x"87",x"cb",x"c1",x"02"),
   288 => (x"ff",x"c0",x"1e",x"c0"),
   289 => (x"49",x"fa",x"c1",x"f0"),
   290 => (x"c4",x"87",x"da",x"f6"),
   291 => (x"9b",x"4b",x"70",x"86"),
   292 => (x"87",x"ed",x"c0",x"05"),
   293 => (x"1e",x"c2",x"cd",x"1e"),
   294 => (x"c3",x"87",x"e1",x"ef"),
   295 => (x"4b",x"6d",x"7d",x"ff"),
   296 => (x"1e",x"ce",x"cd",x"1e"),
   297 => (x"d0",x"87",x"d5",x"ef"),
   298 => (x"7d",x"ff",x"c3",x"86"),
   299 => (x"73",x"7d",x"7d",x"7d"),
   300 => (x"99",x"c0",x"c1",x"49"),
   301 => (x"c1",x"87",x"c5",x"02"),
   302 => (x"87",x"e8",x"c0",x"48"),
   303 => (x"e3",x"c0",x"48",x"c0"),
   304 => (x"cd",x"1e",x"73",x"87"),
   305 => (x"f3",x"ee",x"1e",x"dc"),
   306 => (x"c2",x"86",x"c8",x"87"),
   307 => (x"87",x"cc",x"05",x"ac"),
   308 => (x"ee",x"1e",x"e8",x"cd"),
   309 => (x"86",x"c4",x"87",x"e6"),
   310 => (x"87",x"c8",x"48",x"c0"),
   311 => (x"fe",x"05",x"8c",x"c1"),
   312 => (x"48",x"c0",x"87",x"d5"),
   313 => (x"0e",x"87",x"f6",x"f4"),
   314 => (x"5d",x"5c",x"5b",x"5e"),
   315 => (x"d0",x"ff",x"1e",x"0e"),
   316 => (x"c0",x"c0",x"c8",x"4d"),
   317 => (x"c4",x"f0",x"c2",x"4b"),
   318 => (x"ce",x"78",x"c1",x"48"),
   319 => (x"e6",x"f2",x"49",x"e0"),
   320 => (x"6d",x"4c",x"c7",x"87"),
   321 => (x"c4",x"98",x"73",x"48"),
   322 => (x"98",x"70",x"58",x"a6"),
   323 => (x"6d",x"87",x"cc",x"02"),
   324 => (x"c4",x"98",x"73",x"48"),
   325 => (x"98",x"70",x"58",x"a6"),
   326 => (x"c2",x"87",x"f4",x"05"),
   327 => (x"87",x"fe",x"f5",x"7d"),
   328 => (x"98",x"73",x"48",x"6d"),
   329 => (x"70",x"58",x"a6",x"c4"),
   330 => (x"87",x"cc",x"02",x"98"),
   331 => (x"98",x"73",x"48",x"6d"),
   332 => (x"70",x"58",x"a6",x"c4"),
   333 => (x"87",x"f4",x"05",x"98"),
   334 => (x"1e",x"c0",x"7d",x"c3"),
   335 => (x"c1",x"d0",x"e5",x"c0"),
   336 => (x"e0",x"f3",x"49",x"c0"),
   337 => (x"c1",x"86",x"c4",x"87"),
   338 => (x"87",x"c1",x"05",x"a8"),
   339 => (x"05",x"ac",x"c2",x"4c"),
   340 => (x"db",x"ce",x"87",x"cb"),
   341 => (x"87",x"cf",x"f1",x"49"),
   342 => (x"d8",x"c1",x"48",x"c0"),
   343 => (x"05",x"8c",x"c1",x"87"),
   344 => (x"fb",x"87",x"e0",x"fe"),
   345 => (x"f0",x"c2",x"87",x"c4"),
   346 => (x"98",x"70",x"58",x"c8"),
   347 => (x"c1",x"87",x"cd",x"05"),
   348 => (x"f0",x"ff",x"c0",x"1e"),
   349 => (x"f2",x"49",x"d0",x"c1"),
   350 => (x"86",x"c4",x"87",x"eb"),
   351 => (x"c3",x"48",x"d4",x"ff"),
   352 => (x"e7",x"c5",x"78",x"ff"),
   353 => (x"cc",x"f0",x"c2",x"87"),
   354 => (x"ce",x"1e",x"70",x"58"),
   355 => (x"eb",x"eb",x"1e",x"e4"),
   356 => (x"6d",x"86",x"c8",x"87"),
   357 => (x"c4",x"98",x"73",x"48"),
   358 => (x"98",x"70",x"58",x"a6"),
   359 => (x"6d",x"87",x"cc",x"02"),
   360 => (x"c4",x"98",x"73",x"48"),
   361 => (x"98",x"70",x"58",x"a6"),
   362 => (x"c2",x"87",x"f4",x"05"),
   363 => (x"48",x"d4",x"ff",x"7d"),
   364 => (x"c1",x"78",x"ff",x"c3"),
   365 => (x"e4",x"f1",x"26",x"48"),
   366 => (x"5b",x"5e",x"0e",x"87"),
   367 => (x"1e",x"0e",x"5d",x"5c"),
   368 => (x"4b",x"c0",x"c0",x"c8"),
   369 => (x"ee",x"c5",x"4c",x"c0"),
   370 => (x"c4",x"4a",x"df",x"cd"),
   371 => (x"d4",x"ff",x"5c",x"a6"),
   372 => (x"7c",x"ff",x"c3",x"4c"),
   373 => (x"fe",x"c3",x"48",x"6c"),
   374 => (x"c0",x"c2",x"05",x"a8"),
   375 => (x"05",x"99",x"71",x"87"),
   376 => (x"ff",x"87",x"e2",x"c0"),
   377 => (x"73",x"48",x"bf",x"d0"),
   378 => (x"58",x"a6",x"c4",x"98"),
   379 => (x"ce",x"02",x"98",x"70"),
   380 => (x"bf",x"d0",x"ff",x"87"),
   381 => (x"c4",x"98",x"73",x"48"),
   382 => (x"98",x"70",x"58",x"a6"),
   383 => (x"ff",x"87",x"f2",x"05"),
   384 => (x"d1",x"c4",x"48",x"d0"),
   385 => (x"48",x"66",x"d4",x"78"),
   386 => (x"06",x"a8",x"b7",x"c0"),
   387 => (x"c3",x"87",x"e0",x"c0"),
   388 => (x"4a",x"6c",x"7c",x"ff"),
   389 => (x"c7",x"02",x"99",x"71"),
   390 => (x"97",x"0a",x"71",x"87"),
   391 => (x"81",x"c1",x"0a",x"7a"),
   392 => (x"c1",x"48",x"66",x"d4"),
   393 => (x"58",x"a6",x"d8",x"88"),
   394 => (x"01",x"a8",x"b7",x"c0"),
   395 => (x"c3",x"87",x"e0",x"ff"),
   396 => (x"71",x"7c",x"7c",x"ff"),
   397 => (x"e1",x"c0",x"05",x"99"),
   398 => (x"bf",x"d0",x"ff",x"87"),
   399 => (x"c4",x"98",x"73",x"48"),
   400 => (x"98",x"70",x"58",x"a6"),
   401 => (x"ff",x"87",x"ce",x"02"),
   402 => (x"73",x"48",x"bf",x"d0"),
   403 => (x"58",x"a6",x"c4",x"98"),
   404 => (x"f2",x"05",x"98",x"70"),
   405 => (x"48",x"d0",x"ff",x"87"),
   406 => (x"4a",x"c1",x"78",x"d0"),
   407 => (x"05",x"8a",x"c1",x"7e"),
   408 => (x"6e",x"87",x"ee",x"fd"),
   409 => (x"f4",x"ee",x"26",x"48"),
   410 => (x"5b",x"5e",x"0e",x"87"),
   411 => (x"71",x"1e",x"0e",x"5c"),
   412 => (x"c0",x"c0",x"c8",x"4a"),
   413 => (x"ff",x"4c",x"c0",x"4b"),
   414 => (x"ff",x"c3",x"48",x"d4"),
   415 => (x"bf",x"d0",x"ff",x"78"),
   416 => (x"c4",x"98",x"73",x"48"),
   417 => (x"98",x"70",x"58",x"a6"),
   418 => (x"ff",x"87",x"ce",x"02"),
   419 => (x"73",x"48",x"bf",x"d0"),
   420 => (x"58",x"a6",x"c4",x"98"),
   421 => (x"f2",x"05",x"98",x"70"),
   422 => (x"48",x"d0",x"ff",x"87"),
   423 => (x"ff",x"78",x"c3",x"c4"),
   424 => (x"ff",x"c3",x"48",x"d4"),
   425 => (x"c0",x"1e",x"72",x"78"),
   426 => (x"d1",x"c1",x"f0",x"ff"),
   427 => (x"87",x"f5",x"ed",x"49"),
   428 => (x"98",x"70",x"86",x"c4"),
   429 => (x"87",x"ee",x"c0",x"05"),
   430 => (x"d4",x"1e",x"c0",x"c8"),
   431 => (x"f8",x"fb",x"49",x"66"),
   432 => (x"70",x"86",x"c4",x"87"),
   433 => (x"bf",x"d0",x"ff",x"4c"),
   434 => (x"c4",x"98",x"73",x"48"),
   435 => (x"98",x"70",x"58",x"a6"),
   436 => (x"ff",x"87",x"ce",x"02"),
   437 => (x"73",x"48",x"bf",x"d0"),
   438 => (x"58",x"a6",x"c4",x"98"),
   439 => (x"f2",x"05",x"98",x"70"),
   440 => (x"48",x"d0",x"ff",x"87"),
   441 => (x"48",x"74",x"78",x"c2"),
   442 => (x"87",x"f3",x"ec",x"26"),
   443 => (x"5c",x"5b",x"5e",x"0e"),
   444 => (x"c0",x"1e",x"0e",x"5d"),
   445 => (x"f0",x"ff",x"c0",x"1e"),
   446 => (x"ec",x"49",x"c9",x"c1"),
   447 => (x"1e",x"d2",x"87",x"e7"),
   448 => (x"49",x"d2",x"f0",x"c2"),
   449 => (x"c8",x"87",x"f2",x"fa"),
   450 => (x"c1",x"4d",x"c0",x"86"),
   451 => (x"ad",x"b7",x"d2",x"85"),
   452 => (x"c2",x"87",x"f8",x"04"),
   453 => (x"bf",x"97",x"d2",x"f0"),
   454 => (x"99",x"c0",x"c3",x"49"),
   455 => (x"05",x"a9",x"c0",x"c1"),
   456 => (x"c2",x"87",x"e7",x"c0"),
   457 => (x"bf",x"97",x"d9",x"f0"),
   458 => (x"c2",x"31",x"d0",x"49"),
   459 => (x"bf",x"97",x"da",x"f0"),
   460 => (x"72",x"32",x"c8",x"4a"),
   461 => (x"db",x"f0",x"c2",x"b1"),
   462 => (x"b1",x"4a",x"bf",x"97"),
   463 => (x"ff",x"cf",x"4d",x"71"),
   464 => (x"c1",x"9d",x"ff",x"ff"),
   465 => (x"c2",x"35",x"ca",x"85"),
   466 => (x"f0",x"c2",x"87",x"de"),
   467 => (x"4b",x"bf",x"97",x"db"),
   468 => (x"9b",x"c6",x"33",x"c1"),
   469 => (x"97",x"dc",x"f0",x"c2"),
   470 => (x"b7",x"c7",x"49",x"bf"),
   471 => (x"c2",x"b3",x"71",x"29"),
   472 => (x"bf",x"97",x"d7",x"f0"),
   473 => (x"98",x"cf",x"48",x"49"),
   474 => (x"c2",x"58",x"a6",x"c4"),
   475 => (x"bf",x"97",x"d8",x"f0"),
   476 => (x"ca",x"9c",x"c3",x"4c"),
   477 => (x"d9",x"f0",x"c2",x"34"),
   478 => (x"c2",x"49",x"bf",x"97"),
   479 => (x"c2",x"b4",x"71",x"31"),
   480 => (x"bf",x"97",x"da",x"f0"),
   481 => (x"99",x"c0",x"c3",x"49"),
   482 => (x"71",x"29",x"b7",x"c6"),
   483 => (x"70",x"1e",x"74",x"b4"),
   484 => (x"cf",x"1e",x"73",x"1e"),
   485 => (x"e3",x"e3",x"1e",x"c6"),
   486 => (x"c1",x"83",x"c2",x"87"),
   487 => (x"70",x"30",x"73",x"48"),
   488 => (x"f3",x"cf",x"1e",x"4b"),
   489 => (x"87",x"d4",x"e3",x"1e"),
   490 => (x"66",x"d8",x"48",x"c1"),
   491 => (x"58",x"a6",x"dc",x"30"),
   492 => (x"4d",x"49",x"a4",x"c1"),
   493 => (x"1e",x"70",x"95",x"73"),
   494 => (x"fc",x"cf",x"1e",x"75"),
   495 => (x"87",x"fc",x"e2",x"1e"),
   496 => (x"6e",x"86",x"e4",x"c0"),
   497 => (x"b7",x"c0",x"c8",x"48"),
   498 => (x"87",x"d2",x"06",x"a8"),
   499 => (x"48",x"6e",x"35",x"c1"),
   500 => (x"c4",x"28",x"b7",x"c1"),
   501 => (x"c0",x"c8",x"58",x"a6"),
   502 => (x"ff",x"01",x"a8",x"b7"),
   503 => (x"1e",x"75",x"87",x"ee"),
   504 => (x"e2",x"1e",x"d2",x"d0"),
   505 => (x"86",x"c8",x"87",x"d6"),
   506 => (x"e8",x"26",x"48",x"75"),
   507 => (x"5e",x"0e",x"87",x"ef"),
   508 => (x"71",x"0e",x"5c",x"5b"),
   509 => (x"d0",x"4c",x"c0",x"4b"),
   510 => (x"b7",x"c0",x"48",x"66"),
   511 => (x"e3",x"c0",x"06",x"a8"),
   512 => (x"cc",x"4a",x"13",x"87"),
   513 => (x"49",x"bf",x"97",x"66"),
   514 => (x"c1",x"48",x"66",x"cc"),
   515 => (x"58",x"a6",x"d0",x"80"),
   516 => (x"02",x"aa",x"b7",x"71"),
   517 => (x"48",x"c1",x"87",x"c4"),
   518 => (x"84",x"c1",x"87",x"cc"),
   519 => (x"ac",x"b7",x"66",x"d0"),
   520 => (x"87",x"dd",x"ff",x"04"),
   521 => (x"87",x"c2",x"48",x"c0"),
   522 => (x"4c",x"26",x"4d",x"26"),
   523 => (x"4f",x"26",x"4b",x"26"),
   524 => (x"5c",x"5b",x"5e",x"0e"),
   525 => (x"f8",x"c2",x"0e",x"5d"),
   526 => (x"78",x"c0",x"48",x"f8"),
   527 => (x"49",x"dd",x"ef",x"c0"),
   528 => (x"c2",x"87",x"e4",x"e5"),
   529 => (x"c0",x"1e",x"f0",x"f0"),
   530 => (x"87",x"dd",x"f8",x"49"),
   531 => (x"98",x"70",x"86",x"c4"),
   532 => (x"c0",x"87",x"cc",x"05"),
   533 => (x"e5",x"49",x"c9",x"ec"),
   534 => (x"48",x"c0",x"87",x"cd"),
   535 => (x"c0",x"87",x"e7",x"ca"),
   536 => (x"e5",x"49",x"ea",x"ef"),
   537 => (x"4b",x"c0",x"87",x"c1"),
   538 => (x"48",x"f0",x"fd",x"c2"),
   539 => (x"1e",x"c8",x"78",x"c1"),
   540 => (x"1e",x"c1",x"f0",x"c0"),
   541 => (x"49",x"e6",x"f1",x"c2"),
   542 => (x"c8",x"87",x"f3",x"fd"),
   543 => (x"05",x"98",x"70",x"86"),
   544 => (x"fd",x"c2",x"87",x"c6"),
   545 => (x"78",x"c0",x"48",x"f0"),
   546 => (x"f0",x"c0",x"1e",x"c8"),
   547 => (x"f2",x"c2",x"1e",x"ca"),
   548 => (x"d9",x"fd",x"49",x"c2"),
   549 => (x"70",x"86",x"c8",x"87"),
   550 => (x"87",x"c6",x"05",x"98"),
   551 => (x"48",x"f0",x"fd",x"c2"),
   552 => (x"fd",x"c2",x"78",x"c0"),
   553 => (x"c0",x"1e",x"bf",x"f0"),
   554 => (x"ff",x"1e",x"d3",x"f0"),
   555 => (x"c8",x"87",x"cd",x"df"),
   556 => (x"f0",x"fd",x"c2",x"86"),
   557 => (x"f7",x"c1",x"02",x"bf"),
   558 => (x"ee",x"f8",x"c2",x"87"),
   559 => (x"1e",x"49",x"bf",x"9f"),
   560 => (x"49",x"ee",x"f8",x"c2"),
   561 => (x"a0",x"c2",x"f8",x"48"),
   562 => (x"d0",x"1e",x"71",x"89"),
   563 => (x"1e",x"c0",x"c8",x"1e"),
   564 => (x"1e",x"fb",x"ec",x"c0"),
   565 => (x"87",x"e4",x"de",x"ff"),
   566 => (x"f7",x"c2",x"86",x"d4"),
   567 => (x"c2",x"4b",x"bf",x"f6"),
   568 => (x"bf",x"9f",x"ee",x"f8"),
   569 => (x"ea",x"d6",x"c5",x"4a"),
   570 => (x"c8",x"c0",x"05",x"aa"),
   571 => (x"f6",x"f7",x"c2",x"87"),
   572 => (x"d4",x"c0",x"4b",x"bf"),
   573 => (x"d5",x"e9",x"ca",x"87"),
   574 => (x"cc",x"c0",x"02",x"aa"),
   575 => (x"dd",x"ec",x"c0",x"87"),
   576 => (x"87",x"e3",x"e2",x"49"),
   577 => (x"fd",x"c7",x"48",x"c0"),
   578 => (x"c0",x"1e",x"73",x"87"),
   579 => (x"ff",x"1e",x"f8",x"ed"),
   580 => (x"c2",x"87",x"e9",x"dd"),
   581 => (x"73",x"1e",x"f0",x"f0"),
   582 => (x"87",x"cd",x"f5",x"49"),
   583 => (x"98",x"70",x"86",x"cc"),
   584 => (x"87",x"c5",x"c0",x"05"),
   585 => (x"dd",x"c7",x"48",x"c0"),
   586 => (x"d0",x"ee",x"c0",x"87"),
   587 => (x"87",x"f7",x"e1",x"49"),
   588 => (x"1e",x"e6",x"f0",x"c0"),
   589 => (x"87",x"c4",x"dd",x"ff"),
   590 => (x"f0",x"c0",x"1e",x"c8"),
   591 => (x"f2",x"c2",x"1e",x"fe"),
   592 => (x"e9",x"fa",x"49",x"c2"),
   593 => (x"70",x"86",x"cc",x"87"),
   594 => (x"c9",x"c0",x"05",x"98"),
   595 => (x"f8",x"f8",x"c2",x"87"),
   596 => (x"c0",x"78",x"c1",x"48"),
   597 => (x"1e",x"c8",x"87",x"e4"),
   598 => (x"1e",x"c7",x"f1",x"c0"),
   599 => (x"49",x"e6",x"f1",x"c2"),
   600 => (x"c8",x"87",x"cb",x"fa"),
   601 => (x"02",x"98",x"70",x"86"),
   602 => (x"c0",x"87",x"cf",x"c0"),
   603 => (x"ff",x"1e",x"f7",x"ee"),
   604 => (x"c4",x"87",x"c9",x"dc"),
   605 => (x"c6",x"48",x"c0",x"86"),
   606 => (x"f8",x"c2",x"87",x"cc"),
   607 => (x"49",x"bf",x"97",x"ee"),
   608 => (x"05",x"a9",x"d5",x"c1"),
   609 => (x"c2",x"87",x"cd",x"c0"),
   610 => (x"bf",x"97",x"ef",x"f8"),
   611 => (x"a9",x"ea",x"c2",x"49"),
   612 => (x"87",x"c5",x"c0",x"02"),
   613 => (x"ed",x"c5",x"48",x"c0"),
   614 => (x"f0",x"f0",x"c2",x"87"),
   615 => (x"c3",x"4c",x"bf",x"97"),
   616 => (x"c0",x"02",x"ac",x"e9"),
   617 => (x"eb",x"c3",x"87",x"cc"),
   618 => (x"c5",x"c0",x"02",x"ac"),
   619 => (x"c5",x"48",x"c0",x"87"),
   620 => (x"f0",x"c2",x"87",x"d4"),
   621 => (x"49",x"bf",x"97",x"fb"),
   622 => (x"cc",x"c0",x"05",x"99"),
   623 => (x"fc",x"f0",x"c2",x"87"),
   624 => (x"c2",x"49",x"bf",x"97"),
   625 => (x"c5",x"c0",x"02",x"a9"),
   626 => (x"c4",x"48",x"c0",x"87"),
   627 => (x"f0",x"c2",x"87",x"f8"),
   628 => (x"48",x"bf",x"97",x"fd"),
   629 => (x"58",x"f4",x"f8",x"c2"),
   630 => (x"c1",x"4a",x"49",x"70"),
   631 => (x"f8",x"f8",x"c2",x"8a"),
   632 => (x"71",x"1e",x"72",x"5a"),
   633 => (x"d0",x"f1",x"c0",x"1e"),
   634 => (x"cf",x"da",x"ff",x"1e"),
   635 => (x"c2",x"86",x"cc",x"87"),
   636 => (x"bf",x"97",x"fe",x"f0"),
   637 => (x"c2",x"81",x"73",x"49"),
   638 => (x"bf",x"97",x"ff",x"f0"),
   639 => (x"35",x"c8",x"4d",x"4a"),
   640 => (x"fd",x"c2",x"85",x"71"),
   641 => (x"f1",x"c2",x"5d",x"d0"),
   642 => (x"48",x"bf",x"97",x"c0"),
   643 => (x"58",x"e4",x"fd",x"c2"),
   644 => (x"bf",x"f8",x"f8",x"c2"),
   645 => (x"87",x"dc",x"c2",x"02"),
   646 => (x"ef",x"c0",x"1e",x"c8"),
   647 => (x"f2",x"c2",x"1e",x"d4"),
   648 => (x"c9",x"f7",x"49",x"c2"),
   649 => (x"70",x"86",x"c8",x"87"),
   650 => (x"c5",x"c0",x"02",x"98"),
   651 => (x"c3",x"48",x"c0",x"87"),
   652 => (x"f8",x"c2",x"87",x"d4"),
   653 => (x"48",x"4a",x"bf",x"f0"),
   654 => (x"f9",x"c2",x"30",x"c4"),
   655 => (x"fd",x"c2",x"58",x"c0"),
   656 => (x"f1",x"c2",x"5a",x"e0"),
   657 => (x"49",x"bf",x"97",x"d5"),
   658 => (x"f1",x"c2",x"31",x"c8"),
   659 => (x"4b",x"bf",x"97",x"d4"),
   660 => (x"f1",x"c2",x"49",x"a1"),
   661 => (x"4b",x"bf",x"97",x"d6"),
   662 => (x"a1",x"73",x"33",x"d0"),
   663 => (x"d7",x"f1",x"c2",x"49"),
   664 => (x"d8",x"4b",x"bf",x"97"),
   665 => (x"49",x"a1",x"73",x"33"),
   666 => (x"59",x"e8",x"fd",x"c2"),
   667 => (x"bf",x"e0",x"fd",x"c2"),
   668 => (x"cc",x"fd",x"c2",x"91"),
   669 => (x"fd",x"c2",x"81",x"bf"),
   670 => (x"f1",x"c2",x"59",x"d4"),
   671 => (x"4b",x"bf",x"97",x"dd"),
   672 => (x"f1",x"c2",x"33",x"c8"),
   673 => (x"4c",x"bf",x"97",x"dc"),
   674 => (x"f1",x"c2",x"4b",x"a3"),
   675 => (x"4c",x"bf",x"97",x"de"),
   676 => (x"a3",x"74",x"34",x"d0"),
   677 => (x"df",x"f1",x"c2",x"4b"),
   678 => (x"cf",x"4c",x"bf",x"97"),
   679 => (x"74",x"34",x"d8",x"9c"),
   680 => (x"fd",x"c2",x"4b",x"a3"),
   681 => (x"8b",x"c2",x"5b",x"d8"),
   682 => (x"fd",x"c2",x"92",x"73"),
   683 => (x"a1",x"72",x"48",x"d8"),
   684 => (x"87",x"cb",x"c1",x"78"),
   685 => (x"97",x"c2",x"f1",x"c2"),
   686 => (x"31",x"c8",x"49",x"bf"),
   687 => (x"97",x"c1",x"f1",x"c2"),
   688 => (x"49",x"a1",x"4a",x"bf"),
   689 => (x"59",x"c0",x"f9",x"c2"),
   690 => (x"ff",x"c7",x"31",x"c5"),
   691 => (x"c2",x"29",x"c9",x"81"),
   692 => (x"c2",x"59",x"e0",x"fd"),
   693 => (x"bf",x"97",x"c7",x"f1"),
   694 => (x"c2",x"32",x"c8",x"4a"),
   695 => (x"bf",x"97",x"c6",x"f1"),
   696 => (x"c2",x"4a",x"a2",x"4b"),
   697 => (x"c2",x"5a",x"e8",x"fd"),
   698 => (x"92",x"bf",x"e0",x"fd"),
   699 => (x"fd",x"c2",x"82",x"75"),
   700 => (x"fd",x"c2",x"5a",x"dc"),
   701 => (x"78",x"c0",x"48",x"d4"),
   702 => (x"48",x"d0",x"fd",x"c2"),
   703 => (x"c0",x"78",x"a1",x"72"),
   704 => (x"87",x"e3",x"cd",x"49"),
   705 => (x"df",x"f4",x"48",x"c1"),
   706 => (x"61",x"65",x"52",x"87"),
   707 => (x"66",x"6f",x"20",x"64"),
   708 => (x"52",x"42",x"4d",x"20"),
   709 => (x"69",x"61",x"66",x"20"),
   710 => (x"0a",x"64",x"65",x"6c"),
   711 => (x"20",x"6f",x"4e",x"00"),
   712 => (x"74",x"72",x"61",x"70"),
   713 => (x"6f",x"69",x"74",x"69"),
   714 => (x"69",x"73",x"20",x"6e"),
   715 => (x"74",x"61",x"6e",x"67"),
   716 => (x"20",x"65",x"72",x"75"),
   717 => (x"6e",x"75",x"6f",x"66"),
   718 => (x"4d",x"00",x"0a",x"64"),
   719 => (x"69",x"73",x"52",x"42"),
   720 => (x"20",x"3a",x"65",x"7a"),
   721 => (x"20",x"2c",x"64",x"25"),
   722 => (x"74",x"72",x"61",x"70"),
   723 => (x"6f",x"69",x"74",x"69"),
   724 => (x"7a",x"69",x"73",x"6e"),
   725 => (x"25",x"20",x"3a",x"65"),
   726 => (x"6f",x"20",x"2c",x"64"),
   727 => (x"65",x"73",x"66",x"66"),
   728 => (x"66",x"6f",x"20",x"74"),
   729 => (x"67",x"69",x"73",x"20"),
   730 => (x"64",x"25",x"20",x"3a"),
   731 => (x"69",x"73",x"20",x"2c"),
   732 => (x"78",x"30",x"20",x"67"),
   733 => (x"00",x"0a",x"78",x"25"),
   734 => (x"64",x"61",x"65",x"52"),
   735 => (x"20",x"67",x"6e",x"69"),
   736 => (x"74",x"6f",x"6f",x"62"),
   737 => (x"63",x"65",x"73",x"20"),
   738 => (x"20",x"72",x"6f",x"74"),
   739 => (x"00",x"0a",x"64",x"25"),
   740 => (x"64",x"61",x"65",x"52"),
   741 => (x"6f",x"6f",x"62",x"20"),
   742 => (x"65",x"73",x"20",x"74"),
   743 => (x"72",x"6f",x"74",x"63"),
   744 => (x"6f",x"72",x"66",x"20"),
   745 => (x"69",x"66",x"20",x"6d"),
   746 => (x"20",x"74",x"73",x"72"),
   747 => (x"74",x"72",x"61",x"70"),
   748 => (x"6f",x"69",x"74",x"69"),
   749 => (x"55",x"00",x"0a",x"6e"),
   750 => (x"70",x"75",x"73",x"6e"),
   751 => (x"74",x"72",x"6f",x"70"),
   752 => (x"70",x"20",x"64",x"65"),
   753 => (x"69",x"74",x"72",x"61"),
   754 => (x"6e",x"6f",x"69",x"74"),
   755 => (x"70",x"79",x"74",x"20"),
   756 => (x"00",x"0d",x"21",x"65"),
   757 => (x"33",x"54",x"41",x"46"),
   758 => (x"20",x"20",x"20",x"32"),
   759 => (x"61",x"65",x"52",x"00"),
   760 => (x"67",x"6e",x"69",x"64"),
   761 => (x"52",x"42",x"4d",x"20"),
   762 => (x"42",x"4d",x"00",x"0a"),
   763 => (x"75",x"73",x"20",x"52"),
   764 => (x"73",x"65",x"63",x"63"),
   765 => (x"6c",x"75",x"66",x"73"),
   766 => (x"72",x"20",x"79",x"6c"),
   767 => (x"0a",x"64",x"61",x"65"),
   768 => (x"54",x"41",x"46",x"00"),
   769 => (x"20",x"20",x"36",x"31"),
   770 => (x"41",x"46",x"00",x"20"),
   771 => (x"20",x"32",x"33",x"54"),
   772 => (x"50",x"00",x"20",x"20"),
   773 => (x"69",x"74",x"72",x"61"),
   774 => (x"6e",x"6f",x"69",x"74"),
   775 => (x"6e",x"75",x"6f",x"63"),
   776 => (x"64",x"25",x"20",x"74"),
   777 => (x"75",x"48",x"00",x"0a"),
   778 => (x"6e",x"69",x"74",x"6e"),
   779 => (x"6f",x"66",x"20",x"67"),
   780 => (x"69",x"66",x"20",x"72"),
   781 => (x"79",x"73",x"65",x"6c"),
   782 => (x"6d",x"65",x"74",x"73"),
   783 => (x"41",x"46",x"00",x"0a"),
   784 => (x"20",x"32",x"33",x"54"),
   785 => (x"46",x"00",x"20",x"20"),
   786 => (x"36",x"31",x"54",x"41"),
   787 => (x"00",x"20",x"20",x"20"),
   788 => (x"73",x"75",x"6c",x"43"),
   789 => (x"20",x"72",x"65",x"74"),
   790 => (x"65",x"7a",x"69",x"73"),
   791 => (x"64",x"25",x"20",x"3a"),
   792 => (x"6c",x"43",x"20",x"2c"),
   793 => (x"65",x"74",x"73",x"75"),
   794 => (x"61",x"6d",x"20",x"72"),
   795 => (x"20",x"2c",x"6b",x"73"),
   796 => (x"00",x"0a",x"64",x"25"),
   797 => (x"6e",x"65",x"70",x"4f"),
   798 => (x"66",x"20",x"64",x"65"),
   799 => (x"2c",x"65",x"6c",x"69"),
   800 => (x"61",x"6f",x"6c",x"20"),
   801 => (x"67",x"6e",x"69",x"64"),
   802 => (x"0a",x"2e",x"2e",x"2e"),
   803 => (x"6e",x"61",x"43",x"00"),
   804 => (x"6f",x"20",x"74",x"27"),
   805 => (x"20",x"6e",x"65",x"70"),
   806 => (x"00",x"0a",x"73",x"25"),
   807 => (x"5c",x"5b",x"5e",x"0e"),
   808 => (x"4a",x"71",x"0e",x"5d"),
   809 => (x"bf",x"f8",x"f8",x"c2"),
   810 => (x"72",x"87",x"cc",x"02"),
   811 => (x"2b",x"b7",x"c7",x"4b"),
   812 => (x"ff",x"c1",x"4d",x"72"),
   813 => (x"72",x"87",x"ca",x"9d"),
   814 => (x"2b",x"b7",x"c8",x"4b"),
   815 => (x"ff",x"c3",x"4d",x"72"),
   816 => (x"f0",x"f0",x"c2",x"9d"),
   817 => (x"cc",x"fd",x"c2",x"1e"),
   818 => (x"81",x"73",x"49",x"bf"),
   819 => (x"87",x"d9",x"e6",x"71"),
   820 => (x"98",x"70",x"86",x"c4"),
   821 => (x"c0",x"87",x"c5",x"05"),
   822 => (x"87",x"e6",x"c0",x"48"),
   823 => (x"bf",x"f8",x"f8",x"c2"),
   824 => (x"75",x"87",x"d2",x"02"),
   825 => (x"c2",x"91",x"c4",x"49"),
   826 => (x"69",x"81",x"f0",x"f0"),
   827 => (x"ff",x"ff",x"cf",x"4c"),
   828 => (x"cb",x"9c",x"ff",x"ff"),
   829 => (x"c2",x"49",x"75",x"87"),
   830 => (x"f0",x"f0",x"c2",x"91"),
   831 => (x"4c",x"69",x"9f",x"81"),
   832 => (x"e3",x"ec",x"48",x"74"),
   833 => (x"5b",x"5e",x"0e",x"87"),
   834 => (x"f4",x"0e",x"5d",x"5c"),
   835 => (x"c0",x"4c",x"71",x"86"),
   836 => (x"e8",x"fd",x"c2",x"4b"),
   837 => (x"a6",x"c4",x"7e",x"bf"),
   838 => (x"ec",x"fd",x"c2",x"48"),
   839 => (x"a6",x"c8",x"78",x"bf"),
   840 => (x"c2",x"78",x"c0",x"48"),
   841 => (x"48",x"bf",x"fc",x"f8"),
   842 => (x"c2",x"06",x"a8",x"c0"),
   843 => (x"66",x"c8",x"87",x"e3"),
   844 => (x"05",x"99",x"cf",x"49"),
   845 => (x"f0",x"c2",x"87",x"d8"),
   846 => (x"66",x"c8",x"1e",x"f0"),
   847 => (x"80",x"c1",x"48",x"49"),
   848 => (x"e4",x"58",x"a6",x"cc"),
   849 => (x"86",x"c4",x"87",x"e3"),
   850 => (x"4b",x"f0",x"f0",x"c2"),
   851 => (x"e0",x"c0",x"87",x"c3"),
   852 => (x"4a",x"6b",x"97",x"83"),
   853 => (x"e7",x"c1",x"02",x"9a"),
   854 => (x"aa",x"e5",x"c3",x"87"),
   855 => (x"87",x"e0",x"c1",x"02"),
   856 => (x"97",x"49",x"a3",x"cb"),
   857 => (x"99",x"d8",x"49",x"69"),
   858 => (x"87",x"d4",x"c1",x"05"),
   859 => (x"d0",x"ff",x"49",x"73"),
   860 => (x"1e",x"cb",x"87",x"f5"),
   861 => (x"1e",x"66",x"e0",x"c0"),
   862 => (x"f1",x"e9",x"49",x"73"),
   863 => (x"70",x"86",x"c8",x"87"),
   864 => (x"fb",x"c0",x"05",x"98"),
   865 => (x"4a",x"a3",x"dc",x"87"),
   866 => (x"6a",x"49",x"a4",x"c4"),
   867 => (x"49",x"a3",x"da",x"79"),
   868 => (x"9f",x"4d",x"a4",x"c8"),
   869 => (x"c2",x"7d",x"48",x"69"),
   870 => (x"02",x"bf",x"f8",x"f8"),
   871 => (x"a3",x"d4",x"87",x"d3"),
   872 => (x"49",x"69",x"9f",x"49"),
   873 => (x"99",x"ff",x"ff",x"c0"),
   874 => (x"30",x"d0",x"48",x"71"),
   875 => (x"c2",x"58",x"a6",x"c4"),
   876 => (x"6e",x"7e",x"c0",x"87"),
   877 => (x"70",x"80",x"6d",x"48"),
   878 => (x"c1",x"7c",x"c0",x"7d"),
   879 => (x"87",x"c5",x"c1",x"48"),
   880 => (x"c1",x"48",x"66",x"c8"),
   881 => (x"58",x"a6",x"cc",x"80"),
   882 => (x"bf",x"fc",x"f8",x"c2"),
   883 => (x"dd",x"fd",x"04",x"a8"),
   884 => (x"f8",x"f8",x"c2",x"87"),
   885 => (x"ea",x"c0",x"02",x"bf"),
   886 => (x"fa",x"49",x"6e",x"87"),
   887 => (x"a6",x"c4",x"87",x"fe"),
   888 => (x"cf",x"49",x"70",x"58"),
   889 => (x"f8",x"ff",x"ff",x"ff"),
   890 => (x"d6",x"02",x"a9",x"99"),
   891 => (x"c2",x"49",x"70",x"87"),
   892 => (x"f0",x"f8",x"c2",x"89"),
   893 => (x"fd",x"c2",x"91",x"bf"),
   894 => (x"71",x"48",x"bf",x"d0"),
   895 => (x"58",x"a6",x"c8",x"80"),
   896 => (x"c0",x"87",x"db",x"fc"),
   897 => (x"e8",x"8e",x"f4",x"48"),
   898 => (x"73",x"1e",x"87",x"de"),
   899 => (x"6a",x"4a",x"71",x"1e"),
   900 => (x"71",x"81",x"c1",x"49"),
   901 => (x"f4",x"f8",x"c2",x"7a"),
   902 => (x"cb",x"05",x"99",x"bf"),
   903 => (x"4b",x"a2",x"c8",x"87"),
   904 => (x"f7",x"f9",x"49",x"6b"),
   905 => (x"7b",x"49",x"70",x"87"),
   906 => (x"ff",x"e7",x"48",x"c1"),
   907 => (x"1e",x"73",x"1e",x"87"),
   908 => (x"fd",x"c2",x"4b",x"71"),
   909 => (x"c8",x"49",x"bf",x"d0"),
   910 => (x"4a",x"6a",x"4a",x"a3"),
   911 => (x"f8",x"c2",x"8a",x"c2"),
   912 => (x"72",x"92",x"bf",x"f0"),
   913 => (x"f8",x"c2",x"49",x"a1"),
   914 => (x"6b",x"4a",x"bf",x"f4"),
   915 => (x"49",x"a1",x"72",x"9a"),
   916 => (x"71",x"1e",x"66",x"c8"),
   917 => (x"c4",x"87",x"d2",x"e0"),
   918 => (x"05",x"98",x"70",x"86"),
   919 => (x"48",x"c0",x"87",x"c4"),
   920 => (x"48",x"c1",x"87",x"c2"),
   921 => (x"0e",x"87",x"c5",x"e7"),
   922 => (x"0e",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"c0",x"4a",x"71"),
   924 => (x"c0",x"02",x"9a",x"72"),
   925 => (x"a2",x"da",x"87",x"e0"),
   926 => (x"4b",x"69",x"9f",x"49"),
   927 => (x"bf",x"f8",x"f8",x"c2"),
   928 => (x"d4",x"87",x"cf",x"02"),
   929 => (x"69",x"9f",x"49",x"a2"),
   930 => (x"ff",x"c0",x"4c",x"49"),
   931 => (x"34",x"d0",x"9c",x"ff"),
   932 => (x"4c",x"c0",x"87",x"c2"),
   933 => (x"9b",x"73",x"b3",x"74"),
   934 => (x"4a",x"87",x"df",x"02"),
   935 => (x"f8",x"c2",x"8a",x"c2"),
   936 => (x"92",x"49",x"bf",x"f0"),
   937 => (x"bf",x"d0",x"fd",x"c2"),
   938 => (x"c2",x"80",x"72",x"48"),
   939 => (x"71",x"58",x"f0",x"fd"),
   940 => (x"c2",x"30",x"c4",x"48"),
   941 => (x"c0",x"58",x"c0",x"f9"),
   942 => (x"fd",x"c2",x"87",x"e9"),
   943 => (x"c2",x"4b",x"bf",x"d4"),
   944 => (x"c2",x"48",x"ec",x"fd"),
   945 => (x"78",x"bf",x"d8",x"fd"),
   946 => (x"bf",x"f8",x"f8",x"c2"),
   947 => (x"c2",x"87",x"c9",x"02"),
   948 => (x"49",x"bf",x"f0",x"f8"),
   949 => (x"87",x"c7",x"31",x"c4"),
   950 => (x"bf",x"dc",x"fd",x"c2"),
   951 => (x"c2",x"31",x"c4",x"49"),
   952 => (x"c2",x"59",x"c0",x"f9"),
   953 => (x"e5",x"5b",x"ec",x"fd"),
   954 => (x"5e",x"0e",x"87",x"c0"),
   955 => (x"0e",x"5d",x"5c",x"5b"),
   956 => (x"9a",x"4a",x"71",x"1e"),
   957 => (x"c2",x"87",x"de",x"02"),
   958 => (x"c0",x"48",x"ec",x"f0"),
   959 => (x"e4",x"f0",x"c2",x"78"),
   960 => (x"ec",x"fd",x"c2",x"48"),
   961 => (x"f0",x"c2",x"78",x"bf"),
   962 => (x"fd",x"c2",x"48",x"e8"),
   963 => (x"c1",x"78",x"bf",x"e8"),
   964 => (x"c0",x"48",x"e2",x"c2"),
   965 => (x"fc",x"f8",x"c2",x"78"),
   966 => (x"f0",x"c2",x"49",x"bf"),
   967 => (x"71",x"4a",x"bf",x"ec"),
   968 => (x"fe",x"c3",x"03",x"aa"),
   969 => (x"cf",x"49",x"72",x"87"),
   970 => (x"e1",x"c0",x"05",x"99"),
   971 => (x"f0",x"f0",x"c2",x"87"),
   972 => (x"e4",x"f0",x"c2",x"1e"),
   973 => (x"f0",x"c2",x"49",x"bf"),
   974 => (x"a1",x"c1",x"48",x"e4"),
   975 => (x"dc",x"ff",x"71",x"78"),
   976 => (x"86",x"c4",x"87",x"e7"),
   977 => (x"48",x"de",x"c2",x"c1"),
   978 => (x"78",x"f0",x"f0",x"c2"),
   979 => (x"c2",x"c1",x"87",x"cc"),
   980 => (x"c0",x"48",x"bf",x"de"),
   981 => (x"c2",x"c1",x"80",x"e0"),
   982 => (x"f0",x"c2",x"58",x"e2"),
   983 => (x"c1",x"48",x"bf",x"ec"),
   984 => (x"f0",x"f0",x"c2",x"80"),
   985 => (x"de",x"c2",x"c1",x"58"),
   986 => (x"a3",x"cb",x"4b",x"bf"),
   987 => (x"cf",x"4c",x"11",x"49"),
   988 => (x"dd",x"c1",x"05",x"ac"),
   989 => (x"10",x"9e",x"27",x"87"),
   990 => (x"97",x"bf",x"00",x"00"),
   991 => (x"99",x"df",x"49",x"bf"),
   992 => (x"91",x"cd",x"89",x"c1"),
   993 => (x"81",x"c0",x"f9",x"c2"),
   994 => (x"12",x"4a",x"a3",x"c1"),
   995 => (x"4a",x"a3",x"c3",x"51"),
   996 => (x"a3",x"c5",x"51",x"12"),
   997 => (x"c7",x"51",x"12",x"4a"),
   998 => (x"51",x"12",x"4a",x"a3"),
   999 => (x"12",x"4a",x"a3",x"c9"),
  1000 => (x"4a",x"a3",x"ce",x"51"),
  1001 => (x"a3",x"d0",x"51",x"12"),
  1002 => (x"d2",x"51",x"12",x"4a"),
  1003 => (x"51",x"12",x"4a",x"a3"),
  1004 => (x"12",x"4a",x"a3",x"d4"),
  1005 => (x"4a",x"a3",x"d6",x"51"),
  1006 => (x"a3",x"d8",x"51",x"12"),
  1007 => (x"dc",x"51",x"12",x"4a"),
  1008 => (x"51",x"12",x"4a",x"a3"),
  1009 => (x"12",x"4a",x"a3",x"de"),
  1010 => (x"e2",x"c2",x"c1",x"51"),
  1011 => (x"c1",x"78",x"c1",x"48"),
  1012 => (x"49",x"74",x"87",x"c1"),
  1013 => (x"c0",x"05",x"99",x"c8"),
  1014 => (x"49",x"74",x"87",x"f3"),
  1015 => (x"d0",x"05",x"99",x"d0"),
  1016 => (x"02",x"66",x"d4",x"87"),
  1017 => (x"73",x"87",x"ca",x"c0"),
  1018 => (x"0f",x"66",x"d4",x"49"),
  1019 => (x"dc",x"02",x"98",x"70"),
  1020 => (x"e2",x"c2",x"c1",x"87"),
  1021 => (x"c6",x"c0",x"05",x"bf"),
  1022 => (x"c0",x"f9",x"c2",x"87"),
  1023 => (x"c1",x"50",x"c0",x"48"),
  1024 => (x"c0",x"48",x"e2",x"c2"),
  1025 => (x"de",x"c2",x"c1",x"78"),
  1026 => (x"cc",x"c2",x"48",x"bf"),
  1027 => (x"e2",x"c2",x"c1",x"87"),
  1028 => (x"c2",x"78",x"c0",x"48"),
  1029 => (x"49",x"bf",x"fc",x"f8"),
  1030 => (x"bf",x"ec",x"f0",x"c2"),
  1031 => (x"04",x"aa",x"71",x"4a"),
  1032 => (x"c2",x"87",x"c2",x"fc"),
  1033 => (x"05",x"bf",x"ec",x"fd"),
  1034 => (x"c2",x"87",x"c8",x"c0"),
  1035 => (x"02",x"bf",x"f8",x"f8"),
  1036 => (x"c2",x"87",x"e4",x"c1"),
  1037 => (x"49",x"bf",x"e8",x"f0"),
  1038 => (x"c2",x"87",x"e1",x"f1"),
  1039 => (x"70",x"58",x"ec",x"f0"),
  1040 => (x"f8",x"f8",x"c2",x"4d"),
  1041 => (x"d7",x"c0",x"02",x"bf"),
  1042 => (x"cf",x"49",x"75",x"87"),
  1043 => (x"f8",x"ff",x"ff",x"ff"),
  1044 => (x"c0",x"02",x"a9",x"99"),
  1045 => (x"4c",x"c0",x"87",x"c5"),
  1046 => (x"c1",x"87",x"d9",x"c0"),
  1047 => (x"87",x"d4",x"c0",x"4c"),
  1048 => (x"ff",x"cf",x"49",x"75"),
  1049 => (x"02",x"a9",x"99",x"f8"),
  1050 => (x"c0",x"87",x"c5",x"c0"),
  1051 => (x"87",x"c2",x"c0",x"7e"),
  1052 => (x"4c",x"6e",x"7e",x"c1"),
  1053 => (x"c0",x"05",x"9c",x"74"),
  1054 => (x"49",x"75",x"87",x"dd"),
  1055 => (x"f8",x"c2",x"89",x"c2"),
  1056 => (x"c2",x"91",x"bf",x"f0"),
  1057 => (x"48",x"bf",x"d0",x"fd"),
  1058 => (x"f0",x"c2",x"80",x"71"),
  1059 => (x"f0",x"c2",x"58",x"e8"),
  1060 => (x"78",x"c0",x"48",x"ec"),
  1061 => (x"c0",x"87",x"fe",x"f9"),
  1062 => (x"de",x"ff",x"26",x"48"),
  1063 => (x"00",x"00",x"87",x"ca"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"ff",x"1e",x"00",x"00"),
  1066 => (x"ff",x"c3",x"48",x"d4"),
  1067 => (x"99",x"49",x"68",x"78"),
  1068 => (x"c0",x"87",x"c6",x"02"),
  1069 => (x"ee",x"05",x"a9",x"fb"),
  1070 => (x"26",x"48",x"71",x"87"),
  1071 => (x"5b",x"5e",x"0e",x"4f"),
  1072 => (x"4a",x"71",x"0e",x"5c"),
  1073 => (x"d4",x"ff",x"4b",x"c0"),
  1074 => (x"78",x"ff",x"c3",x"48"),
  1075 => (x"02",x"99",x"49",x"68"),
  1076 => (x"c0",x"87",x"c1",x"c1"),
  1077 => (x"c0",x"02",x"a9",x"ec"),
  1078 => (x"fb",x"c0",x"87",x"fa"),
  1079 => (x"f3",x"c0",x"02",x"a9"),
  1080 => (x"b7",x"66",x"cc",x"87"),
  1081 => (x"87",x"cc",x"03",x"ab"),
  1082 => (x"c7",x"02",x"66",x"d0"),
  1083 => (x"97",x"09",x"72",x"87"),
  1084 => (x"82",x"c1",x"09",x"79"),
  1085 => (x"c2",x"02",x"99",x"71"),
  1086 => (x"ff",x"83",x"c1",x"87"),
  1087 => (x"ff",x"c3",x"48",x"d4"),
  1088 => (x"99",x"49",x"68",x"78"),
  1089 => (x"c0",x"87",x"cd",x"02"),
  1090 => (x"c7",x"02",x"a9",x"ec"),
  1091 => (x"a9",x"fb",x"c0",x"87"),
  1092 => (x"87",x"cd",x"ff",x"05"),
  1093 => (x"c3",x"02",x"66",x"d0"),
  1094 => (x"7a",x"97",x"c0",x"87"),
  1095 => (x"05",x"a9",x"fb",x"c0"),
  1096 => (x"4c",x"73",x"87",x"c7"),
  1097 => (x"c2",x"8c",x"0c",x"c0"),
  1098 => (x"74",x"4c",x"73",x"87"),
  1099 => (x"26",x"87",x"c2",x"48"),
  1100 => (x"26",x"4c",x"26",x"4d"),
  1101 => (x"1e",x"4f",x"26",x"4b"),
  1102 => (x"c3",x"48",x"d4",x"ff"),
  1103 => (x"49",x"68",x"78",x"ff"),
  1104 => (x"a9",x"b7",x"f0",x"c0"),
  1105 => (x"c0",x"87",x"ca",x"04"),
  1106 => (x"01",x"a9",x"b7",x"f9"),
  1107 => (x"f0",x"c0",x"87",x"c3"),
  1108 => (x"b7",x"c1",x"c1",x"89"),
  1109 => (x"87",x"ca",x"04",x"a9"),
  1110 => (x"a9",x"b7",x"c6",x"c1"),
  1111 => (x"c0",x"87",x"c3",x"01"),
  1112 => (x"48",x"71",x"89",x"f7"),
  1113 => (x"5e",x"0e",x"4f",x"26"),
  1114 => (x"0e",x"5d",x"5c",x"5b"),
  1115 => (x"4c",x"71",x"86",x"f4"),
  1116 => (x"c0",x"4b",x"d4",x"ff"),
  1117 => (x"ff",x"c3",x"7e",x"4d"),
  1118 => (x"bf",x"d0",x"ff",x"7b"),
  1119 => (x"c0",x"c0",x"c8",x"48"),
  1120 => (x"58",x"a6",x"c8",x"98"),
  1121 => (x"d0",x"02",x"98",x"70"),
  1122 => (x"bf",x"d0",x"ff",x"87"),
  1123 => (x"c0",x"c0",x"c8",x"48"),
  1124 => (x"58",x"a6",x"c8",x"98"),
  1125 => (x"f0",x"05",x"98",x"70"),
  1126 => (x"48",x"d0",x"ff",x"87"),
  1127 => (x"d4",x"78",x"e1",x"c0"),
  1128 => (x"87",x"c2",x"fc",x"7b"),
  1129 => (x"02",x"99",x"49",x"70"),
  1130 => (x"c3",x"87",x"c7",x"c1"),
  1131 => (x"a6",x"c8",x"7b",x"ff"),
  1132 => (x"c8",x"78",x"6b",x"48"),
  1133 => (x"fb",x"c0",x"48",x"66"),
  1134 => (x"87",x"c8",x"02",x"a8"),
  1135 => (x"bf",x"c8",x"fe",x"c2"),
  1136 => (x"87",x"ee",x"c0",x"02"),
  1137 => (x"99",x"71",x"4d",x"c1"),
  1138 => (x"87",x"e6",x"c0",x"02"),
  1139 => (x"02",x"a9",x"fb",x"c0"),
  1140 => (x"d1",x"fb",x"87",x"c3"),
  1141 => (x"7b",x"ff",x"c3",x"87"),
  1142 => (x"c6",x"c1",x"49",x"6b"),
  1143 => (x"87",x"cc",x"05",x"a9"),
  1144 => (x"7b",x"7b",x"ff",x"c3"),
  1145 => (x"6b",x"48",x"a6",x"c8"),
  1146 => (x"4d",x"49",x"c0",x"78"),
  1147 => (x"ff",x"05",x"99",x"71"),
  1148 => (x"9d",x"75",x"87",x"da"),
  1149 => (x"87",x"de",x"c1",x"05"),
  1150 => (x"6b",x"7b",x"ff",x"c3"),
  1151 => (x"7b",x"ff",x"c3",x"4a"),
  1152 => (x"6b",x"48",x"a6",x"c4"),
  1153 => (x"c1",x"48",x"6e",x"78"),
  1154 => (x"58",x"a6",x"c4",x"80"),
  1155 => (x"97",x"49",x"a4",x"c8"),
  1156 => (x"66",x"c8",x"49",x"69"),
  1157 => (x"87",x"da",x"05",x"a9"),
  1158 => (x"97",x"49",x"a4",x"c9"),
  1159 => (x"05",x"aa",x"49",x"69"),
  1160 => (x"a4",x"ca",x"87",x"d0"),
  1161 => (x"49",x"69",x"97",x"49"),
  1162 => (x"05",x"a9",x"66",x"c4"),
  1163 => (x"4d",x"c1",x"87",x"c4"),
  1164 => (x"66",x"c8",x"87",x"d6"),
  1165 => (x"a8",x"ec",x"c0",x"48"),
  1166 => (x"c8",x"87",x"c9",x"02"),
  1167 => (x"fb",x"c0",x"48",x"66"),
  1168 => (x"87",x"c4",x"05",x"a8"),
  1169 => (x"4d",x"c1",x"7e",x"c0"),
  1170 => (x"c8",x"7b",x"ff",x"c3"),
  1171 => (x"78",x"6b",x"48",x"a6"),
  1172 => (x"fe",x"02",x"9d",x"75"),
  1173 => (x"d0",x"ff",x"87",x"e2"),
  1174 => (x"c0",x"c8",x"48",x"bf"),
  1175 => (x"a6",x"c8",x"98",x"c0"),
  1176 => (x"02",x"98",x"70",x"58"),
  1177 => (x"d0",x"ff",x"87",x"d0"),
  1178 => (x"c0",x"c8",x"48",x"bf"),
  1179 => (x"a6",x"c8",x"98",x"c0"),
  1180 => (x"05",x"98",x"70",x"58"),
  1181 => (x"d0",x"ff",x"87",x"f0"),
  1182 => (x"78",x"e0",x"c0",x"48"),
  1183 => (x"8e",x"f4",x"48",x"6e"),
  1184 => (x"0e",x"87",x"ec",x"fa"),
  1185 => (x"5d",x"5c",x"5b",x"5e"),
  1186 => (x"d0",x"ff",x"1e",x"0e"),
  1187 => (x"c0",x"c0",x"c8",x"4b"),
  1188 => (x"d0",x"fe",x"c2",x"4a"),
  1189 => (x"48",x"6b",x"4d",x"bf"),
  1190 => (x"a6",x"c4",x"98",x"72"),
  1191 => (x"02",x"98",x"70",x"58"),
  1192 => (x"48",x"6b",x"87",x"cc"),
  1193 => (x"a6",x"c4",x"98",x"72"),
  1194 => (x"05",x"98",x"70",x"58"),
  1195 => (x"7b",x"c5",x"87",x"f4"),
  1196 => (x"c1",x"48",x"d4",x"ff"),
  1197 => (x"78",x"c3",x"78",x"d3"),
  1198 => (x"98",x"72",x"48",x"6b"),
  1199 => (x"70",x"58",x"a6",x"c4"),
  1200 => (x"87",x"cc",x"02",x"98"),
  1201 => (x"98",x"72",x"48",x"6b"),
  1202 => (x"70",x"58",x"a6",x"c4"),
  1203 => (x"87",x"f4",x"05",x"98"),
  1204 => (x"48",x"6b",x"7b",x"c4"),
  1205 => (x"a6",x"c4",x"98",x"72"),
  1206 => (x"02",x"98",x"70",x"58"),
  1207 => (x"48",x"6b",x"87",x"cc"),
  1208 => (x"a6",x"c4",x"98",x"72"),
  1209 => (x"05",x"98",x"70",x"58"),
  1210 => (x"d1",x"c4",x"87",x"f4"),
  1211 => (x"02",x"9d",x"75",x"7b"),
  1212 => (x"c8",x"87",x"f2",x"c0"),
  1213 => (x"04",x"ad",x"b7",x"c0"),
  1214 => (x"8d",x"4a",x"87",x"c4"),
  1215 => (x"4a",x"75",x"87",x"c4"),
  1216 => (x"49",x"72",x"4d",x"c0"),
  1217 => (x"99",x"71",x"8a",x"c1"),
  1218 => (x"ff",x"87",x"ce",x"02"),
  1219 => (x"78",x"c0",x"48",x"d4"),
  1220 => (x"8a",x"c1",x"49",x"72"),
  1221 => (x"f2",x"05",x"99",x"71"),
  1222 => (x"48",x"d4",x"ff",x"87"),
  1223 => (x"75",x"78",x"78",x"c0"),
  1224 => (x"ce",x"ff",x"05",x"9d"),
  1225 => (x"c0",x"c0",x"c8",x"87"),
  1226 => (x"72",x"48",x"6b",x"4a"),
  1227 => (x"58",x"a6",x"c4",x"98"),
  1228 => (x"cc",x"02",x"98",x"70"),
  1229 => (x"72",x"48",x"6b",x"87"),
  1230 => (x"58",x"a6",x"c4",x"98"),
  1231 => (x"f4",x"05",x"98",x"70"),
  1232 => (x"6b",x"7b",x"d0",x"87"),
  1233 => (x"c4",x"98",x"72",x"48"),
  1234 => (x"98",x"70",x"58",x"a6"),
  1235 => (x"6b",x"87",x"cc",x"02"),
  1236 => (x"c4",x"98",x"72",x"48"),
  1237 => (x"98",x"70",x"58",x"a6"),
  1238 => (x"c5",x"87",x"f4",x"05"),
  1239 => (x"48",x"d4",x"ff",x"7b"),
  1240 => (x"c0",x"78",x"d3",x"c1"),
  1241 => (x"72",x"48",x"6b",x"78"),
  1242 => (x"58",x"a6",x"c4",x"98"),
  1243 => (x"cc",x"02",x"98",x"70"),
  1244 => (x"72",x"48",x"6b",x"87"),
  1245 => (x"58",x"a6",x"c4",x"98"),
  1246 => (x"f4",x"05",x"98",x"70"),
  1247 => (x"26",x"7b",x"c4",x"87"),
  1248 => (x"0e",x"87",x"ec",x"f6"),
  1249 => (x"5d",x"5c",x"5b",x"5e"),
  1250 => (x"71",x"86",x"f4",x"0e"),
  1251 => (x"4c",x"d0",x"ff",x"4d"),
  1252 => (x"4b",x"c0",x"c0",x"c8"),
  1253 => (x"fe",x"c2",x"1e",x"75"),
  1254 => (x"e8",x"e5",x"49",x"cc"),
  1255 => (x"70",x"86",x"c4",x"87"),
  1256 => (x"c4",x"c6",x"02",x"98"),
  1257 => (x"d0",x"fe",x"c2",x"87"),
  1258 => (x"49",x"75",x"7e",x"bf"),
  1259 => (x"c8",x"87",x"f7",x"f6"),
  1260 => (x"1e",x"70",x"58",x"a6"),
  1261 => (x"1e",x"49",x"a5",x"c8"),
  1262 => (x"1e",x"c0",x"d5",x"c1"),
  1263 => (x"87",x"fc",x"f2",x"fe"),
  1264 => (x"48",x"6c",x"86",x"cc"),
  1265 => (x"a6",x"cc",x"98",x"73"),
  1266 => (x"02",x"98",x"70",x"58"),
  1267 => (x"48",x"6c",x"87",x"cc"),
  1268 => (x"a6",x"cc",x"98",x"73"),
  1269 => (x"05",x"98",x"70",x"58"),
  1270 => (x"7c",x"c5",x"87",x"f4"),
  1271 => (x"c1",x"48",x"d4",x"ff"),
  1272 => (x"fe",x"c2",x"78",x"d5"),
  1273 => (x"c1",x"49",x"bf",x"c8"),
  1274 => (x"4a",x"66",x"c4",x"81"),
  1275 => (x"32",x"c6",x"8a",x"c1"),
  1276 => (x"b0",x"71",x"48",x"72"),
  1277 => (x"78",x"08",x"d4",x"ff"),
  1278 => (x"98",x"73",x"48",x"6c"),
  1279 => (x"70",x"58",x"a6",x"cc"),
  1280 => (x"87",x"cc",x"02",x"98"),
  1281 => (x"98",x"73",x"48",x"6c"),
  1282 => (x"70",x"58",x"a6",x"c8"),
  1283 => (x"87",x"f4",x"05",x"98"),
  1284 => (x"d4",x"ff",x"7c",x"c4"),
  1285 => (x"78",x"ff",x"c3",x"48"),
  1286 => (x"98",x"73",x"48",x"6c"),
  1287 => (x"70",x"58",x"a6",x"c8"),
  1288 => (x"87",x"cc",x"02",x"98"),
  1289 => (x"98",x"73",x"48",x"6c"),
  1290 => (x"70",x"58",x"a6",x"c8"),
  1291 => (x"87",x"f4",x"05",x"98"),
  1292 => (x"d4",x"ff",x"7c",x"c5"),
  1293 => (x"78",x"d3",x"c1",x"48"),
  1294 => (x"48",x"6c",x"78",x"c1"),
  1295 => (x"a6",x"c8",x"98",x"73"),
  1296 => (x"02",x"98",x"70",x"58"),
  1297 => (x"48",x"6c",x"87",x"cc"),
  1298 => (x"a6",x"c8",x"98",x"73"),
  1299 => (x"05",x"98",x"70",x"58"),
  1300 => (x"7c",x"c4",x"87",x"f4"),
  1301 => (x"d0",x"c2",x"02",x"6e"),
  1302 => (x"f0",x"f0",x"c2",x"87"),
  1303 => (x"fe",x"c2",x"1e",x"4d"),
  1304 => (x"c8",x"e7",x"49",x"cc"),
  1305 => (x"70",x"86",x"c4",x"87"),
  1306 => (x"87",x"c5",x"05",x"98"),
  1307 => (x"ca",x"c3",x"48",x"c0"),
  1308 => (x"c8",x"48",x"6e",x"87"),
  1309 => (x"04",x"a8",x"b7",x"c0"),
  1310 => (x"6e",x"4a",x"87",x"cb"),
  1311 => (x"88",x"c0",x"c8",x"48"),
  1312 => (x"c4",x"58",x"a6",x"c4"),
  1313 => (x"c0",x"4a",x"6e",x"87"),
  1314 => (x"73",x"48",x"6c",x"7e"),
  1315 => (x"58",x"a6",x"c8",x"98"),
  1316 => (x"cc",x"02",x"98",x"70"),
  1317 => (x"73",x"48",x"6c",x"87"),
  1318 => (x"58",x"a6",x"c8",x"98"),
  1319 => (x"f4",x"05",x"98",x"70"),
  1320 => (x"ff",x"7c",x"cd",x"87"),
  1321 => (x"d4",x"c1",x"48",x"d4"),
  1322 => (x"c1",x"49",x"72",x"78"),
  1323 => (x"02",x"99",x"71",x"8a"),
  1324 => (x"48",x"15",x"87",x"d0"),
  1325 => (x"78",x"08",x"d4",x"ff"),
  1326 => (x"8a",x"c1",x"49",x"72"),
  1327 => (x"ff",x"05",x"99",x"71"),
  1328 => (x"48",x"6c",x"87",x"f0"),
  1329 => (x"a6",x"c8",x"98",x"73"),
  1330 => (x"02",x"98",x"70",x"58"),
  1331 => (x"48",x"6c",x"87",x"cd"),
  1332 => (x"a6",x"c8",x"98",x"73"),
  1333 => (x"05",x"98",x"70",x"58"),
  1334 => (x"c4",x"87",x"f3",x"ff"),
  1335 => (x"cc",x"fe",x"c2",x"7c"),
  1336 => (x"87",x"e6",x"e4",x"49"),
  1337 => (x"f0",x"fd",x"05",x"6e"),
  1338 => (x"73",x"48",x"6c",x"87"),
  1339 => (x"58",x"a6",x"c4",x"98"),
  1340 => (x"cd",x"02",x"98",x"70"),
  1341 => (x"73",x"48",x"6c",x"87"),
  1342 => (x"58",x"a6",x"c4",x"98"),
  1343 => (x"ff",x"05",x"98",x"70"),
  1344 => (x"7c",x"c5",x"87",x"f3"),
  1345 => (x"c1",x"48",x"d4",x"ff"),
  1346 => (x"78",x"c0",x"78",x"d3"),
  1347 => (x"98",x"73",x"48",x"6c"),
  1348 => (x"70",x"58",x"a6",x"c4"),
  1349 => (x"87",x"cd",x"02",x"98"),
  1350 => (x"98",x"73",x"48",x"6c"),
  1351 => (x"70",x"58",x"a6",x"c4"),
  1352 => (x"f3",x"ff",x"05",x"98"),
  1353 => (x"d0",x"7c",x"c4",x"87"),
  1354 => (x"c1",x"1e",x"75",x"87"),
  1355 => (x"fe",x"1e",x"e6",x"d5"),
  1356 => (x"c8",x"87",x"c9",x"ed"),
  1357 => (x"c2",x"48",x"c0",x"86"),
  1358 => (x"f4",x"48",x"c1",x"87"),
  1359 => (x"87",x"ef",x"ef",x"8e"),
  1360 => (x"6e",x"65",x"70",x"4f"),
  1361 => (x"66",x"20",x"64",x"65"),
  1362 => (x"2c",x"65",x"6c",x"69"),
  1363 => (x"61",x"6f",x"6c",x"20"),
  1364 => (x"67",x"6e",x"69",x"64"),
  1365 => (x"2c",x"73",x"25",x"20"),
  1366 => (x"64",x"69",x"28",x"20"),
  1367 => (x"64",x"25",x"20",x"78"),
  1368 => (x"2e",x"2e",x"2e",x"29"),
  1369 => (x"61",x"43",x"00",x"0a"),
  1370 => (x"20",x"74",x"27",x"6e"),
  1371 => (x"6e",x"65",x"70",x"6f"),
  1372 => (x"0a",x"73",x"25",x"20"),
  1373 => (x"6f",x"6f",x"4c",x"00"),
  1374 => (x"67",x"6e",x"69",x"6b"),
  1375 => (x"72",x"6f",x"66",x"20"),
  1376 => (x"6c",x"69",x"66",x"20"),
  1377 => (x"64",x"25",x"20",x"65"),
  1378 => (x"69",x"46",x"00",x"0a"),
  1379 => (x"25",x"20",x"65",x"6c"),
  1380 => (x"53",x"00",x"0a",x"73"),
  1381 => (x"63",x"65",x"6c",x"65"),
  1382 => (x"20",x"64",x"65",x"74"),
  1383 => (x"6d",x"6f",x"72",x"66"),
  1384 => (x"20",x"64",x"25",x"20"),
  1385 => (x"64",x"25",x"20",x"2b"),
  1386 => (x"69",x"6c",x"00",x"0a"),
  1387 => (x"6f",x"72",x"74",x"73"),
  1388 => (x"6b",x"73",x"20",x"6d"),
  1389 => (x"69",x"70",x"70",x"69"),
  1390 => (x"25",x"20",x"67",x"6e"),
  1391 => (x"64",x"20",x"2c",x"64"),
  1392 => (x"6e",x"65",x"72",x"69"),
  1393 => (x"65",x"69",x"72",x"74"),
  1394 => (x"64",x"25",x"20",x"73"),
  1395 => (x"80",x"00",x"0a",x"20"),
  1396 => (x"63",x"61",x"42",x"20"),
  1397 => (x"75",x"73",x"00",x"6b"),
  1398 => (x"6e",x"65",x"6d",x"62"),
  1399 => (x"61",x"63",x"20",x"75"),
  1400 => (x"61",x"62",x"6c",x"6c"),
  1401 => (x"4c",x"00",x"6b",x"63"),
  1402 => (x"20",x"64",x"61",x"6f"),
  1403 => (x"00",x"20",x"2e",x"2a"),
  1404 => (x"64",x"61",x"6f",x"4c"),
  1405 => (x"00",x"20",x"3a",x"00"),
  1406 => (x"6f",x"63",x"65",x"44"),
  1407 => (x"20",x"64",x"65",x"64"),
  1408 => (x"6f",x"20",x"64",x"25"),
  1409 => (x"6f",x"69",x"74",x"70"),
  1410 => (x"00",x"0a",x"73",x"6e"),
  1411 => (x"65",x"67",x"61",x"50"),
  1412 => (x"0a",x"64",x"25",x"20"),
  1413 => (x"42",x"20",x"80",x"00"),
  1414 => (x"00",x"6b",x"63",x"61"),
  1415 => (x"78",x"45",x"20",x"80"),
  1416 => (x"4e",x"00",x"74",x"69"),
  1417 => (x"20",x"74",x"78",x"65"),
  1418 => (x"72",x"61",x"68",x"63"),
  1419 => (x"0a",x"63",x"25",x"20"),
  1420 => (x"78",x"61",x"4d",x"00"),
  1421 => (x"65",x"67",x"61",x"70"),
  1422 => (x"0a",x"64",x"25",x"20"),
  1423 => (x"4d",x"4f",x"52",x"00"),
  1424 => (x"61",x"6f",x"6c",x"20"),
  1425 => (x"0a",x"64",x"65",x"64"),
  1426 => (x"4d",x"4f",x"52",x"00"),
  1427 => (x"61",x"6f",x"6c",x"20"),
  1428 => (x"61",x"66",x"20",x"64"),
  1429 => (x"64",x"65",x"6c",x"69"),
  1430 => (x"6e",x"49",x"00",x"0a"),
  1431 => (x"61",x"69",x"74",x"69"),
  1432 => (x"69",x"7a",x"69",x"6c"),
  1433 => (x"53",x"20",x"67",x"6e"),
  1434 => (x"61",x"63",x"20",x"44"),
  1435 => (x"00",x"0a",x"64",x"72"),
  1436 => (x"65",x"76",x"61",x"48"),
  1437 => (x"0a",x"44",x"53",x"20"),
  1438 => (x"5b",x"5e",x"0e",x"00"),
  1439 => (x"1e",x"0e",x"5d",x"5c"),
  1440 => (x"4c",x"c0",x"4b",x"71"),
  1441 => (x"d5",x"c1",x"1e",x"73"),
  1442 => (x"e7",x"fe",x"1e",x"f5"),
  1443 => (x"86",x"c8",x"87",x"ee"),
  1444 => (x"ab",x"b7",x"4d",x"c0"),
  1445 => (x"87",x"e9",x"c0",x"04"),
  1446 => (x"1e",x"e6",x"c5",x"c1"),
  1447 => (x"c4",x"02",x"9d",x"75"),
  1448 => (x"c2",x"4a",x"c0",x"87"),
  1449 => (x"72",x"4a",x"c1",x"87"),
  1450 => (x"87",x"fe",x"e0",x"49"),
  1451 => (x"58",x"a6",x"86",x"c4"),
  1452 => (x"05",x"6e",x"84",x"c1"),
  1453 => (x"4c",x"73",x"87",x"c2"),
  1454 => (x"b7",x"73",x"85",x"c1"),
  1455 => (x"d7",x"ff",x"06",x"ac"),
  1456 => (x"26",x"48",x"6e",x"87"),
  1457 => (x"0e",x"87",x"e8",x"e9"),
  1458 => (x"5d",x"5c",x"5b",x"5e"),
  1459 => (x"1e",x"4c",x"71",x"0e"),
  1460 => (x"bf",x"d8",x"fe",x"c2"),
  1461 => (x"d3",x"d6",x"c1",x"1e"),
  1462 => (x"df",x"e6",x"fe",x"1e"),
  1463 => (x"d8",x"fe",x"c2",x"87"),
  1464 => (x"81",x"74",x"49",x"bf"),
  1465 => (x"70",x"87",x"d2",x"fe"),
  1466 => (x"d6",x"c1",x"1e",x"4d"),
  1467 => (x"e6",x"fe",x"1e",x"ca"),
  1468 => (x"86",x"d4",x"87",x"ca"),
  1469 => (x"d3",x"02",x"9d",x"75"),
  1470 => (x"c0",x"f9",x"c2",x"87"),
  1471 => (x"cb",x"4a",x"75",x"4b"),
  1472 => (x"c6",x"eb",x"fe",x"49"),
  1473 => (x"c0",x"f9",x"c2",x"87"),
  1474 => (x"87",x"f7",x"f1",x"49"),
  1475 => (x"49",x"fd",x"fb",x"c1"),
  1476 => (x"87",x"c6",x"c7",x"c1"),
  1477 => (x"87",x"e2",x"c7",x"c1"),
  1478 => (x"1e",x"87",x"d4",x"e8"),
  1479 => (x"4b",x"71",x"1e",x"73"),
  1480 => (x"d8",x"fe",x"c2",x"49"),
  1481 => (x"d0",x"fd",x"81",x"bf"),
  1482 => (x"9a",x"4a",x"70",x"87"),
  1483 => (x"49",x"87",x"c5",x"02"),
  1484 => (x"87",x"f3",x"dc",x"ff"),
  1485 => (x"48",x"d8",x"fe",x"c2"),
  1486 => (x"49",x"73",x"78",x"c0"),
  1487 => (x"e7",x"87",x"e9",x"c1"),
  1488 => (x"73",x"1e",x"87",x"f1"),
  1489 => (x"c4",x"4b",x"71",x"1e"),
  1490 => (x"c1",x"02",x"4a",x"a3"),
  1491 => (x"8a",x"c1",x"87",x"c8"),
  1492 => (x"8a",x"87",x"dc",x"02"),
  1493 => (x"87",x"f1",x"c0",x"02"),
  1494 => (x"c4",x"c1",x"05",x"8a"),
  1495 => (x"d8",x"fe",x"c2",x"87"),
  1496 => (x"fc",x"c0",x"02",x"bf"),
  1497 => (x"88",x"c1",x"48",x"87"),
  1498 => (x"58",x"dc",x"fe",x"c2"),
  1499 => (x"c2",x"87",x"f2",x"c0"),
  1500 => (x"49",x"bf",x"d8",x"fe"),
  1501 => (x"fe",x"c2",x"89",x"d0"),
  1502 => (x"b7",x"c0",x"59",x"dc"),
  1503 => (x"e0",x"c0",x"03",x"a9"),
  1504 => (x"d8",x"fe",x"c2",x"87"),
  1505 => (x"d8",x"78",x"c0",x"48"),
  1506 => (x"d8",x"fe",x"c2",x"87"),
  1507 => (x"80",x"c1",x"48",x"bf"),
  1508 => (x"58",x"dc",x"fe",x"c2"),
  1509 => (x"fe",x"c2",x"87",x"cb"),
  1510 => (x"d0",x"48",x"bf",x"d8"),
  1511 => (x"dc",x"fe",x"c2",x"80"),
  1512 => (x"c3",x"49",x"73",x"58"),
  1513 => (x"87",x"cb",x"e6",x"87"),
  1514 => (x"5c",x"5b",x"5e",x"0e"),
  1515 => (x"86",x"f0",x"0e",x"5d"),
  1516 => (x"c2",x"59",x"a6",x"d0"),
  1517 => (x"c0",x"4d",x"f0",x"f0"),
  1518 => (x"fc",x"f8",x"c2",x"4c"),
  1519 => (x"fe",x"c2",x"1e",x"bf"),
  1520 => (x"c1",x"1e",x"bf",x"d8"),
  1521 => (x"fe",x"1e",x"ea",x"d6"),
  1522 => (x"cc",x"87",x"f1",x"e2"),
  1523 => (x"48",x"a6",x"c4",x"86"),
  1524 => (x"fe",x"c2",x"78",x"c0"),
  1525 => (x"c0",x"48",x"bf",x"d8"),
  1526 => (x"c1",x"06",x"a8",x"b7"),
  1527 => (x"f0",x"c2",x"87",x"c2"),
  1528 => (x"02",x"98",x"48",x"f0"),
  1529 => (x"c1",x"87",x"f9",x"c0"),
  1530 => (x"c8",x"1e",x"e6",x"c5"),
  1531 => (x"87",x"c7",x"02",x"66"),
  1532 => (x"c0",x"48",x"a6",x"c4"),
  1533 => (x"c4",x"87",x"c5",x"78"),
  1534 => (x"78",x"c1",x"48",x"a6"),
  1535 => (x"ff",x"49",x"66",x"c4"),
  1536 => (x"c4",x"87",x"e7",x"db"),
  1537 => (x"c1",x"4d",x"70",x"86"),
  1538 => (x"48",x"66",x"c4",x"84"),
  1539 => (x"a6",x"c8",x"80",x"c1"),
  1540 => (x"d8",x"fe",x"c2",x"58"),
  1541 => (x"03",x"ac",x"b7",x"bf"),
  1542 => (x"9d",x"75",x"87",x"c6"),
  1543 => (x"87",x"c7",x"ff",x"05"),
  1544 => (x"9d",x"75",x"4c",x"c0"),
  1545 => (x"87",x"e5",x"c3",x"02"),
  1546 => (x"1e",x"e6",x"c5",x"c1"),
  1547 => (x"c7",x"02",x"66",x"c8"),
  1548 => (x"48",x"a6",x"cc",x"87"),
  1549 => (x"87",x"c5",x"78",x"c0"),
  1550 => (x"c1",x"48",x"a6",x"cc"),
  1551 => (x"49",x"66",x"cc",x"78"),
  1552 => (x"87",x"e6",x"da",x"ff"),
  1553 => (x"58",x"a6",x"86",x"c4"),
  1554 => (x"ec",x"c2",x"02",x"6e"),
  1555 => (x"81",x"cb",x"49",x"87"),
  1556 => (x"d0",x"49",x"69",x"97"),
  1557 => (x"d9",x"c1",x"02",x"99"),
  1558 => (x"db",x"dc",x"c1",x"87"),
  1559 => (x"cc",x"49",x"74",x"4b"),
  1560 => (x"fd",x"fb",x"c1",x"91"),
  1561 => (x"4a",x"a1",x"c8",x"81"),
  1562 => (x"81",x"c1",x"7a",x"73"),
  1563 => (x"74",x"51",x"ff",x"c3"),
  1564 => (x"c2",x"91",x"de",x"49"),
  1565 => (x"71",x"4d",x"ec",x"fe"),
  1566 => (x"97",x"c1",x"c2",x"85"),
  1567 => (x"49",x"a5",x"c1",x"7d"),
  1568 => (x"c2",x"51",x"e0",x"c0"),
  1569 => (x"bf",x"97",x"c0",x"f9"),
  1570 => (x"c1",x"87",x"d2",x"02"),
  1571 => (x"4b",x"a5",x"c2",x"84"),
  1572 => (x"4a",x"c0",x"f9",x"c2"),
  1573 => (x"e4",x"fe",x"49",x"db"),
  1574 => (x"dc",x"c1",x"87",x"f1"),
  1575 => (x"49",x"a5",x"cd",x"87"),
  1576 => (x"84",x"c1",x"51",x"c0"),
  1577 => (x"6e",x"4b",x"a5",x"c2"),
  1578 => (x"fe",x"49",x"cb",x"4a"),
  1579 => (x"c1",x"87",x"dc",x"e4"),
  1580 => (x"49",x"74",x"87",x"c7"),
  1581 => (x"fb",x"c1",x"91",x"cc"),
  1582 => (x"81",x"c8",x"81",x"fd"),
  1583 => (x"79",x"c7",x"db",x"c1"),
  1584 => (x"97",x"c0",x"f9",x"c2"),
  1585 => (x"87",x"d9",x"02",x"bf"),
  1586 => (x"91",x"de",x"49",x"74"),
  1587 => (x"fe",x"c2",x"84",x"c1"),
  1588 => (x"83",x"71",x"4b",x"ec"),
  1589 => (x"4a",x"c0",x"f9",x"c2"),
  1590 => (x"e3",x"fe",x"49",x"dd"),
  1591 => (x"d8",x"c0",x"87",x"ed"),
  1592 => (x"de",x"4b",x"74",x"87"),
  1593 => (x"ec",x"fe",x"c2",x"93"),
  1594 => (x"49",x"a3",x"cb",x"83"),
  1595 => (x"84",x"c1",x"51",x"c0"),
  1596 => (x"cb",x"4a",x"6e",x"73"),
  1597 => (x"d2",x"e3",x"fe",x"49"),
  1598 => (x"48",x"66",x"c4",x"87"),
  1599 => (x"a6",x"c8",x"80",x"c1"),
  1600 => (x"ac",x"b7",x"c7",x"58"),
  1601 => (x"87",x"c5",x"c0",x"03"),
  1602 => (x"db",x"fc",x"05",x"6e"),
  1603 => (x"ac",x"b7",x"c7",x"87"),
  1604 => (x"87",x"d3",x"c0",x"03"),
  1605 => (x"91",x"de",x"49",x"74"),
  1606 => (x"81",x"ec",x"fe",x"c2"),
  1607 => (x"84",x"c1",x"51",x"c0"),
  1608 => (x"04",x"ac",x"b7",x"c7"),
  1609 => (x"c1",x"87",x"ed",x"ff"),
  1610 => (x"c0",x"48",x"d2",x"fd"),
  1611 => (x"d1",x"fd",x"c1",x"50"),
  1612 => (x"c1",x"50",x"c2",x"48"),
  1613 => (x"c1",x"48",x"d9",x"fd"),
  1614 => (x"c1",x"78",x"e6",x"e5"),
  1615 => (x"c1",x"48",x"d5",x"fd"),
  1616 => (x"c1",x"78",x"cf",x"d7"),
  1617 => (x"c1",x"48",x"e5",x"fd"),
  1618 => (x"cc",x"78",x"c2",x"dd"),
  1619 => (x"fa",x"c0",x"49",x"66"),
  1620 => (x"8e",x"f0",x"87",x"c9"),
  1621 => (x"87",x"d7",x"df",x"ff"),
  1622 => (x"c2",x"4a",x"71",x"1e"),
  1623 => (x"72",x"5a",x"cc",x"fe"),
  1624 => (x"87",x"c4",x"f9",x"49"),
  1625 => (x"73",x"1e",x"4f",x"26"),
  1626 => (x"49",x"4b",x"71",x"1e"),
  1627 => (x"fb",x"c1",x"91",x"cc"),
  1628 => (x"81",x"c1",x"81",x"fd"),
  1629 => (x"fe",x"c2",x"48",x"11"),
  1630 => (x"d7",x"c1",x"58",x"c8"),
  1631 => (x"e0",x"fe",x"49",x"d6"),
  1632 => (x"f0",x"c0",x"87",x"e5"),
  1633 => (x"e1",x"fe",x"49",x"a3"),
  1634 => (x"49",x"c0",x"87",x"d1"),
  1635 => (x"ff",x"87",x"f8",x"d2"),
  1636 => (x"0e",x"87",x"e0",x"de"),
  1637 => (x"5d",x"5c",x"5b",x"5e"),
  1638 => (x"71",x"86",x"f0",x"0e"),
  1639 => (x"91",x"cc",x"49",x"4c"),
  1640 => (x"81",x"fd",x"fb",x"c1"),
  1641 => (x"c4",x"7e",x"a1",x"c3"),
  1642 => (x"fe",x"c2",x"48",x"a6"),
  1643 => (x"6e",x"78",x"bf",x"c0"),
  1644 => (x"c4",x"4a",x"bf",x"97"),
  1645 => (x"2b",x"72",x"4b",x"66"),
  1646 => (x"12",x"4a",x"a1",x"c1"),
  1647 => (x"58",x"a6",x"cc",x"48"),
  1648 => (x"83",x"c1",x"9b",x"70"),
  1649 => (x"69",x"97",x"81",x"c2"),
  1650 => (x"04",x"ab",x"b7",x"49"),
  1651 => (x"4b",x"c0",x"87",x"c2"),
  1652 => (x"4a",x"bf",x"97",x"6e"),
  1653 => (x"72",x"49",x"66",x"c8"),
  1654 => (x"c4",x"b9",x"ff",x"31"),
  1655 => (x"4d",x"73",x"99",x"66"),
  1656 => (x"b5",x"71",x"35",x"72"),
  1657 => (x"5d",x"c4",x"fe",x"c2"),
  1658 => (x"c3",x"48",x"d4",x"ff"),
  1659 => (x"d0",x"ff",x"78",x"ff"),
  1660 => (x"c0",x"c8",x"48",x"bf"),
  1661 => (x"a6",x"d0",x"98",x"c0"),
  1662 => (x"02",x"98",x"70",x"58"),
  1663 => (x"d0",x"ff",x"87",x"d0"),
  1664 => (x"c0",x"c8",x"48",x"bf"),
  1665 => (x"a6",x"c4",x"98",x"c0"),
  1666 => (x"05",x"98",x"70",x"58"),
  1667 => (x"d0",x"ff",x"87",x"f0"),
  1668 => (x"78",x"e1",x"c0",x"48"),
  1669 => (x"de",x"48",x"d4",x"ff"),
  1670 => (x"7d",x"0d",x"70",x"78"),
  1671 => (x"c8",x"48",x"75",x"0d"),
  1672 => (x"d4",x"ff",x"28",x"b7"),
  1673 => (x"48",x"75",x"78",x"08"),
  1674 => (x"ff",x"28",x"b7",x"d0"),
  1675 => (x"75",x"78",x"08",x"d4"),
  1676 => (x"28",x"b7",x"d8",x"48"),
  1677 => (x"78",x"08",x"d4",x"ff"),
  1678 => (x"48",x"bf",x"d0",x"ff"),
  1679 => (x"98",x"c0",x"c0",x"c8"),
  1680 => (x"70",x"58",x"a6",x"c4"),
  1681 => (x"87",x"d0",x"02",x"98"),
  1682 => (x"48",x"bf",x"d0",x"ff"),
  1683 => (x"98",x"c0",x"c0",x"c8"),
  1684 => (x"70",x"58",x"a6",x"c4"),
  1685 => (x"87",x"f0",x"05",x"98"),
  1686 => (x"c0",x"48",x"d0",x"ff"),
  1687 => (x"1e",x"c7",x"78",x"e0"),
  1688 => (x"fb",x"c1",x"1e",x"c0"),
  1689 => (x"fe",x"c2",x"1e",x"fd"),
  1690 => (x"cc",x"49",x"bf",x"c4"),
  1691 => (x"c0",x"49",x"74",x"87"),
  1692 => (x"e4",x"87",x"e8",x"f5"),
  1693 => (x"f6",x"da",x"ff",x"8e"),
  1694 => (x"5b",x"5e",x"0e",x"87"),
  1695 => (x"ff",x"0e",x"5d",x"5c"),
  1696 => (x"a6",x"d8",x"86",x"d8"),
  1697 => (x"48",x"a6",x"c8",x"59"),
  1698 => (x"80",x"c4",x"78",x"c0"),
  1699 => (x"80",x"c4",x"78",x"c0"),
  1700 => (x"d4",x"ff",x"78",x"c0"),
  1701 => (x"78",x"ff",x"c3",x"48"),
  1702 => (x"48",x"bf",x"d0",x"ff"),
  1703 => (x"98",x"c0",x"c0",x"c8"),
  1704 => (x"70",x"58",x"a6",x"c4"),
  1705 => (x"87",x"d0",x"02",x"98"),
  1706 => (x"48",x"bf",x"d0",x"ff"),
  1707 => (x"98",x"c0",x"c0",x"c8"),
  1708 => (x"70",x"58",x"a6",x"c4"),
  1709 => (x"87",x"f0",x"05",x"98"),
  1710 => (x"c0",x"48",x"d0",x"ff"),
  1711 => (x"d4",x"ff",x"78",x"e1"),
  1712 => (x"ff",x"78",x"d4",x"48"),
  1713 => (x"ff",x"87",x"df",x"d7"),
  1714 => (x"ff",x"c3",x"48",x"d4"),
  1715 => (x"1e",x"4d",x"68",x"78"),
  1716 => (x"1e",x"e3",x"d8",x"c1"),
  1717 => (x"87",x"e4",x"d6",x"fe"),
  1718 => (x"fb",x"c0",x"86",x"c8"),
  1719 => (x"c5",x"c1",x"02",x"ad"),
  1720 => (x"66",x"f8",x"c0",x"87"),
  1721 => (x"6a",x"82",x"c4",x"4a"),
  1722 => (x"c1",x"1e",x"72",x"7e"),
  1723 => (x"c4",x"48",x"e7",x"d7"),
  1724 => (x"a1",x"c8",x"49",x"66"),
  1725 => (x"71",x"41",x"20",x"4a"),
  1726 => (x"87",x"f9",x"05",x"aa"),
  1727 => (x"4a",x"26",x"51",x"10"),
  1728 => (x"49",x"66",x"f8",x"c0"),
  1729 => (x"e5",x"c1",x"81",x"c8"),
  1730 => (x"49",x"6a",x"79",x"d8"),
  1731 => (x"0d",x"71",x"81",x"c8"),
  1732 => (x"c1",x"0d",x"7d",x"97"),
  1733 => (x"6a",x"1e",x"d8",x"1e"),
  1734 => (x"ff",x"81",x"c8",x"49"),
  1735 => (x"c8",x"87",x"de",x"d6"),
  1736 => (x"48",x"a6",x"d0",x"86"),
  1737 => (x"9d",x"75",x"78",x"c1"),
  1738 => (x"87",x"e8",x"c9",x"02"),
  1739 => (x"c1",x"48",x"66",x"d0"),
  1740 => (x"a8",x"b7",x"66",x"c0"),
  1741 => (x"87",x"dc",x"c9",x"03"),
  1742 => (x"c3",x"48",x"d4",x"ff"),
  1743 => (x"48",x"68",x"78",x"ff"),
  1744 => (x"c4",x"88",x"c6",x"c1"),
  1745 => (x"98",x"70",x"58",x"a6"),
  1746 => (x"48",x"87",x"db",x"02"),
  1747 => (x"a6",x"c4",x"88",x"c9"),
  1748 => (x"02",x"98",x"70",x"58"),
  1749 => (x"48",x"87",x"eb",x"c3"),
  1750 => (x"a6",x"c4",x"88",x"c1"),
  1751 => (x"02",x"98",x"70",x"58"),
  1752 => (x"c8",x"87",x"c5",x"c1"),
  1753 => (x"66",x"d4",x"87",x"d6"),
  1754 => (x"87",x"f3",x"c0",x"05"),
  1755 => (x"cc",x"49",x"66",x"d0"),
  1756 => (x"66",x"f8",x"c0",x"91"),
  1757 => (x"4a",x"a1",x"c4",x"81"),
  1758 => (x"1e",x"71",x"7e",x"6a"),
  1759 => (x"48",x"f0",x"d7",x"c1"),
  1760 => (x"c4",x"49",x"66",x"c4"),
  1761 => (x"41",x"20",x"4a",x"a1"),
  1762 => (x"f9",x"05",x"aa",x"71"),
  1763 => (x"26",x"51",x"10",x"87"),
  1764 => (x"c1",x"81",x"c8",x"49"),
  1765 => (x"d0",x"79",x"d8",x"e5"),
  1766 => (x"80",x"c1",x"48",x"66"),
  1767 => (x"ff",x"58",x"a6",x"d4"),
  1768 => (x"70",x"87",x"c3",x"d4"),
  1769 => (x"87",x"da",x"c7",x"4d"),
  1770 => (x"87",x"cb",x"d6",x"ff"),
  1771 => (x"70",x"58",x"a6",x"cc"),
  1772 => (x"cc",x"d8",x"c1",x"1e"),
  1773 => (x"c3",x"d3",x"fe",x"1e"),
  1774 => (x"66",x"86",x"c8",x"87"),
  1775 => (x"b7",x"66",x"cc",x"48"),
  1776 => (x"87",x"c6",x"06",x"a8"),
  1777 => (x"c8",x"48",x"a6",x"cc"),
  1778 => (x"d5",x"ff",x"78",x"66"),
  1779 => (x"ec",x"c0",x"87",x"e9"),
  1780 => (x"ed",x"c1",x"05",x"a8"),
  1781 => (x"05",x"66",x"d4",x"87"),
  1782 => (x"d0",x"87",x"de",x"c1"),
  1783 => (x"91",x"cc",x"49",x"66"),
  1784 => (x"81",x"66",x"f8",x"c0"),
  1785 => (x"6a",x"4a",x"a1",x"c4"),
  1786 => (x"4a",x"a1",x"c1",x"4c"),
  1787 => (x"c2",x"52",x"66",x"c8"),
  1788 => (x"81",x"c8",x"79",x"97"),
  1789 => (x"79",x"e6",x"e5",x"c1"),
  1790 => (x"c3",x"48",x"d4",x"ff"),
  1791 => (x"4d",x"68",x"78",x"ff"),
  1792 => (x"e0",x"c0",x"02",x"9d"),
  1793 => (x"ad",x"fb",x"c0",x"87"),
  1794 => (x"74",x"87",x"da",x"02"),
  1795 => (x"0d",x"7d",x"97",x"0d"),
  1796 => (x"d4",x"ff",x"84",x"c1"),
  1797 => (x"78",x"ff",x"c3",x"48"),
  1798 => (x"02",x"9d",x"4d",x"68"),
  1799 => (x"fb",x"c0",x"87",x"c7"),
  1800 => (x"e6",x"ff",x"05",x"ad"),
  1801 => (x"54",x"e0",x"c0",x"87"),
  1802 => (x"c0",x"54",x"c1",x"c2"),
  1803 => (x"66",x"d0",x"7c",x"97"),
  1804 => (x"d4",x"80",x"c1",x"48"),
  1805 => (x"c9",x"c5",x"58",x"a6"),
  1806 => (x"e9",x"d1",x"ff",x"87"),
  1807 => (x"c5",x"4d",x"70",x"87"),
  1808 => (x"66",x"c8",x"87",x"c0"),
  1809 => (x"a8",x"66",x"d4",x"48"),
  1810 => (x"87",x"e7",x"c4",x"05"),
  1811 => (x"c0",x"48",x"a6",x"d8"),
  1812 => (x"e2",x"d3",x"ff",x"78"),
  1813 => (x"a6",x"e0",x"c0",x"87"),
  1814 => (x"da",x"d3",x"ff",x"58"),
  1815 => (x"a6",x"e4",x"c0",x"87"),
  1816 => (x"a8",x"ec",x"c0",x"58"),
  1817 => (x"87",x"ca",x"c0",x"05"),
  1818 => (x"48",x"a6",x"e0",x"c0"),
  1819 => (x"c0",x"78",x"66",x"dc"),
  1820 => (x"d4",x"ff",x"87",x"c6"),
  1821 => (x"78",x"ff",x"c3",x"48"),
  1822 => (x"cc",x"49",x"66",x"d0"),
  1823 => (x"66",x"f8",x"c0",x"91"),
  1824 => (x"c4",x"80",x"71",x"48"),
  1825 => (x"49",x"6e",x"58",x"a6"),
  1826 => (x"66",x"dc",x"81",x"c3"),
  1827 => (x"66",x"e0",x"c0",x"51"),
  1828 => (x"dc",x"81",x"c1",x"49"),
  1829 => (x"48",x"c1",x"89",x"66"),
  1830 => (x"49",x"70",x"30",x"71"),
  1831 => (x"4a",x"6e",x"89",x"c1"),
  1832 => (x"09",x"72",x"82",x"c1"),
  1833 => (x"6e",x"09",x"79",x"97"),
  1834 => (x"6e",x"50",x"c2",x"48"),
  1835 => (x"c1",x"81",x"c8",x"49"),
  1836 => (x"c2",x"79",x"d3",x"e6"),
  1837 => (x"49",x"bf",x"c0",x"fe"),
  1838 => (x"29",x"b7",x"66",x"dc"),
  1839 => (x"48",x"4a",x"6a",x"97"),
  1840 => (x"e8",x"c0",x"98",x"71"),
  1841 => (x"48",x"6e",x"58",x"a6"),
  1842 => (x"a6",x"c8",x"80",x"c4"),
  1843 => (x"bf",x"66",x"c4",x"58"),
  1844 => (x"48",x"66",x"d4",x"4c"),
  1845 => (x"02",x"a8",x"66",x"c8"),
  1846 => (x"dc",x"87",x"c8",x"c0"),
  1847 => (x"78",x"c0",x"48",x"a6"),
  1848 => (x"dc",x"87",x"c5",x"c0"),
  1849 => (x"78",x"c1",x"48",x"a6"),
  1850 => (x"c0",x"1e",x"66",x"dc"),
  1851 => (x"49",x"74",x"1e",x"e0"),
  1852 => (x"87",x"c9",x"cf",x"ff"),
  1853 => (x"4d",x"70",x"86",x"c8"),
  1854 => (x"06",x"ad",x"b7",x"c0"),
  1855 => (x"75",x"87",x"d5",x"c1"),
  1856 => (x"bf",x"66",x"c4",x"84"),
  1857 => (x"81",x"e0",x"c0",x"49"),
  1858 => (x"c1",x"4b",x"89",x"74"),
  1859 => (x"71",x"4a",x"f5",x"d7"),
  1860 => (x"87",x"f7",x"d2",x"fe"),
  1861 => (x"66",x"d8",x"84",x"c2"),
  1862 => (x"dc",x"80",x"c1",x"48"),
  1863 => (x"e4",x"c0",x"58",x"a6"),
  1864 => (x"81",x"c1",x"49",x"66"),
  1865 => (x"c0",x"02",x"a9",x"70"),
  1866 => (x"a6",x"dc",x"87",x"c8"),
  1867 => (x"c0",x"78",x"c0",x"48"),
  1868 => (x"a6",x"dc",x"87",x"c5"),
  1869 => (x"dc",x"78",x"c1",x"48"),
  1870 => (x"66",x"c8",x"1e",x"66"),
  1871 => (x"e0",x"c0",x"49",x"bf"),
  1872 => (x"71",x"89",x"74",x"81"),
  1873 => (x"ff",x"49",x"74",x"1e"),
  1874 => (x"c8",x"87",x"f2",x"cd"),
  1875 => (x"a8",x"b7",x"c0",x"86"),
  1876 => (x"87",x"c2",x"ff",x"01"),
  1877 => (x"c1",x"1e",x"66",x"d8"),
  1878 => (x"fe",x"1e",x"f8",x"d7"),
  1879 => (x"c8",x"87",x"dd",x"cc"),
  1880 => (x"c2",x"49",x"6e",x"86"),
  1881 => (x"51",x"66",x"d8",x"81"),
  1882 => (x"c1",x"48",x"66",x"d0"),
  1883 => (x"58",x"a6",x"d4",x"80"),
  1884 => (x"ff",x"87",x"cf",x"c0"),
  1885 => (x"70",x"87",x"ef",x"cc"),
  1886 => (x"87",x"c6",x"c0",x"4d"),
  1887 => (x"87",x"e6",x"cc",x"ff"),
  1888 => (x"9d",x"75",x"4d",x"70"),
  1889 => (x"87",x"cc",x"c0",x"02"),
  1890 => (x"c1",x"48",x"66",x"d0"),
  1891 => (x"a8",x"b7",x"66",x"c0"),
  1892 => (x"87",x"e4",x"f6",x"04"),
  1893 => (x"c7",x"48",x"66",x"d0"),
  1894 => (x"c0",x"03",x"a8",x"b7"),
  1895 => (x"66",x"d0",x"87",x"e3"),
  1896 => (x"c0",x"91",x"cc",x"49"),
  1897 => (x"c4",x"81",x"66",x"f8"),
  1898 => (x"4a",x"6a",x"4a",x"a1"),
  1899 => (x"81",x"c8",x"52",x"c0"),
  1900 => (x"66",x"d0",x"79",x"c0"),
  1901 => (x"d4",x"80",x"c1",x"48"),
  1902 => (x"b7",x"c7",x"58",x"a6"),
  1903 => (x"dd",x"ff",x"04",x"a8"),
  1904 => (x"02",x"66",x"d4",x"87"),
  1905 => (x"c0",x"87",x"eb",x"c0"),
  1906 => (x"c1",x"49",x"66",x"f8"),
  1907 => (x"f8",x"c0",x"81",x"d4"),
  1908 => (x"d5",x"c1",x"4a",x"66"),
  1909 => (x"c2",x"52",x"c0",x"82"),
  1910 => (x"66",x"f8",x"c0",x"51"),
  1911 => (x"81",x"dc",x"c1",x"49"),
  1912 => (x"79",x"e6",x"e5",x"c1"),
  1913 => (x"49",x"66",x"f8",x"c0"),
  1914 => (x"c1",x"81",x"d8",x"c1"),
  1915 => (x"c0",x"79",x"d5",x"d8"),
  1916 => (x"f8",x"c0",x"87",x"d6"),
  1917 => (x"d8",x"c1",x"49",x"66"),
  1918 => (x"dc",x"d8",x"c1",x"81"),
  1919 => (x"66",x"f8",x"c0",x"79"),
  1920 => (x"81",x"dc",x"c1",x"49"),
  1921 => (x"79",x"fa",x"e3",x"c2"),
  1922 => (x"c1",x"1e",x"66",x"cc"),
  1923 => (x"fe",x"1e",x"f1",x"d8"),
  1924 => (x"c8",x"87",x"e9",x"c9"),
  1925 => (x"bf",x"d0",x"ff",x"86"),
  1926 => (x"c0",x"c0",x"c8",x"48"),
  1927 => (x"58",x"a6",x"c4",x"98"),
  1928 => (x"c0",x"02",x"98",x"70"),
  1929 => (x"d0",x"ff",x"87",x"d1"),
  1930 => (x"c0",x"c8",x"48",x"bf"),
  1931 => (x"a6",x"c4",x"98",x"c0"),
  1932 => (x"05",x"98",x"70",x"58"),
  1933 => (x"ff",x"87",x"ef",x"ff"),
  1934 => (x"e0",x"c0",x"48",x"d0"),
  1935 => (x"48",x"66",x"cc",x"78"),
  1936 => (x"ff",x"8e",x"d8",x"ff"),
  1937 => (x"1e",x"87",x"e8",x"cb"),
  1938 => (x"1e",x"c0",x"1e",x"c7"),
  1939 => (x"1e",x"fd",x"fb",x"c1"),
  1940 => (x"bf",x"c4",x"fe",x"c2"),
  1941 => (x"87",x"e1",x"f0",x"49"),
  1942 => (x"49",x"fd",x"fb",x"c1"),
  1943 => (x"87",x"fa",x"e9",x"c0"),
  1944 => (x"4f",x"26",x"8e",x"f4"),
  1945 => (x"ca",x"1e",x"73",x"1e"),
  1946 => (x"fe",x"c2",x"87",x"f4"),
  1947 => (x"50",x"c0",x"48",x"dc"),
  1948 => (x"c3",x"48",x"d4",x"ff"),
  1949 => (x"d9",x"c1",x"78",x"ff"),
  1950 => (x"cc",x"fe",x"49",x"da"),
  1951 => (x"d9",x"fe",x"87",x"e9"),
  1952 => (x"98",x"70",x"87",x"e5"),
  1953 => (x"fe",x"87",x"cd",x"02"),
  1954 => (x"70",x"87",x"e5",x"e6"),
  1955 => (x"87",x"c4",x"02",x"98"),
  1956 => (x"87",x"c2",x"4b",x"c1"),
  1957 => (x"9b",x"73",x"4b",x"c0"),
  1958 => (x"c1",x"87",x"c8",x"02"),
  1959 => (x"fe",x"49",x"f0",x"d9"),
  1960 => (x"c2",x"87",x"c4",x"cc"),
  1961 => (x"c0",x"48",x"c4",x"fe"),
  1962 => (x"da",x"fe",x"49",x"78"),
  1963 => (x"87",x"da",x"c4",x"87"),
  1964 => (x"c0",x"87",x"ff",x"c9"),
  1965 => (x"c5",x"87",x"d2",x"ea"),
  1966 => (x"87",x"c0",x"ce",x"49"),
  1967 => (x"c4",x"02",x"98",x"70"),
  1968 => (x"fe",x"ce",x"ff",x"87"),
  1969 => (x"49",x"f8",x"c1",x"87"),
  1970 => (x"70",x"87",x"f1",x"cd"),
  1971 => (x"df",x"ff",x"02",x"98"),
  1972 => (x"02",x"9b",x"73",x"87"),
  1973 => (x"fe",x"c2",x"87",x"d8"),
  1974 => (x"d2",x"ff",x"49",x"dc"),
  1975 => (x"98",x"70",x"87",x"e5"),
  1976 => (x"c1",x"87",x"cb",x"02"),
  1977 => (x"fe",x"49",x"fd",x"d8"),
  1978 => (x"ff",x"87",x"fc",x"ca"),
  1979 => (x"d9",x"c1",x"87",x"c2"),
  1980 => (x"ca",x"fe",x"49",x"c9"),
  1981 => (x"f7",x"fe",x"87",x"f1"),
  1982 => (x"f6",x"c8",x"ff",x"87"),
  1983 => (x"00",x"00",x"02",x"87"),
  1984 => (x"00",x"2f",x"ac",x"00"),
  1985 => (x"00",x"16",x"c7",x"00"),
  1986 => (x"00",x"00",x"02",x"00"),
  1987 => (x"00",x"2f",x"ca",x"00"),
  1988 => (x"00",x"16",x"c7",x"00"),
  1989 => (x"00",x"00",x"02",x"00"),
  1990 => (x"00",x"2f",x"e8",x"00"),
  1991 => (x"00",x"16",x"c7",x"00"),
  1992 => (x"00",x"00",x"02",x"00"),
  1993 => (x"00",x"30",x"06",x"00"),
  1994 => (x"00",x"16",x"c7",x"00"),
  1995 => (x"00",x"00",x"02",x"00"),
  1996 => (x"00",x"30",x"24",x"00"),
  1997 => (x"00",x"16",x"c7",x"00"),
  1998 => (x"00",x"00",x"02",x"00"),
  1999 => (x"00",x"30",x"42",x"00"),
  2000 => (x"00",x"16",x"c7",x"00"),
  2001 => (x"00",x"00",x"02",x"00"),
  2002 => (x"00",x"30",x"60",x"00"),
  2003 => (x"00",x"16",x"c7",x"00"),
  2004 => (x"00",x"00",x"02",x"00"),
  2005 => (x"00",x"00",x"00",x"00"),
  2006 => (x"00",x"19",x"66",x"00"),
  2007 => (x"00",x"00",x"00",x"00"),
  2008 => (x"00",x"00",x"00",x"00"),
  2009 => (x"00",x"17",x"42",x"00"),
  2010 => (x"c1",x"1e",x"1e",x"00"),
  2011 => (x"a6",x"c4",x"87",x"d5"),
  2012 => (x"4f",x"26",x"26",x"58"),
  2013 => (x"fe",x"4a",x"71",x"1e"),
  2014 => (x"78",x"c0",x"48",x"f0"),
  2015 => (x"0a",x"7a",x"0a",x"cd"),
  2016 => (x"49",x"ca",x"fe",x"c1"),
  2017 => (x"87",x"df",x"c8",x"fe"),
  2018 => (x"65",x"53",x"4f",x"26"),
  2019 => (x"61",x"68",x"20",x"74"),
  2020 => (x"65",x"6c",x"64",x"6e"),
  2021 => (x"49",x"00",x"0a",x"72"),
  2022 => (x"6e",x"69",x"20",x"6e"),
  2023 => (x"72",x"72",x"65",x"74"),
  2024 => (x"20",x"74",x"70",x"75"),
  2025 => (x"73",x"6e",x"6f",x"63"),
  2026 => (x"63",x"75",x"72",x"74"),
  2027 => (x"0a",x"72",x"6f",x"74"),
  2028 => (x"fe",x"c1",x"1e",x"00"),
  2029 => (x"c7",x"fe",x"49",x"d7"),
  2030 => (x"fd",x"c1",x"87",x"ed"),
  2031 => (x"f3",x"fe",x"49",x"e9"),
  2032 => (x"1e",x"4f",x"26",x"87"),
  2033 => (x"48",x"bf",x"f0",x"fe"),
  2034 => (x"fe",x"1e",x"4f",x"26"),
  2035 => (x"78",x"c1",x"48",x"f0"),
  2036 => (x"fe",x"1e",x"4f",x"26"),
  2037 => (x"78",x"c0",x"48",x"f0"),
  2038 => (x"71",x"1e",x"4f",x"26"),
  2039 => (x"c4",x"7a",x"c0",x"4a"),
  2040 => (x"79",x"c0",x"49",x"a2"),
  2041 => (x"c0",x"49",x"a2",x"c8"),
  2042 => (x"49",x"a2",x"cc",x"79"),
  2043 => (x"4f",x"26",x"79",x"c0"),
  2044 => (x"5c",x"5b",x"5e",x"0e"),
  2045 => (x"71",x"86",x"f8",x"0e"),
  2046 => (x"49",x"a4",x"c8",x"4c"),
  2047 => (x"6b",x"4b",x"a4",x"cc"),
  2048 => (x"c4",x"80",x"c1",x"48"),
  2049 => (x"98",x"cf",x"58",x"a6"),
  2050 => (x"69",x"58",x"a6",x"c8"),
  2051 => (x"a8",x"66",x"c4",x"48"),
  2052 => (x"6b",x"87",x"d4",x"05"),
  2053 => (x"c4",x"80",x"c1",x"48"),
  2054 => (x"98",x"cf",x"58",x"a6"),
  2055 => (x"69",x"58",x"a6",x"c8"),
  2056 => (x"a8",x"66",x"c4",x"48"),
  2057 => (x"fe",x"87",x"ec",x"02"),
  2058 => (x"d0",x"c1",x"87",x"e8"),
  2059 => (x"48",x"6b",x"49",x"a4"),
  2060 => (x"a6",x"c4",x"90",x"c4"),
  2061 => (x"d4",x"81",x"70",x"58"),
  2062 => (x"48",x"6b",x"79",x"66"),
  2063 => (x"a6",x"c8",x"80",x"c1"),
  2064 => (x"70",x"98",x"cf",x"58"),
  2065 => (x"87",x"d2",x"c1",x"7b"),
  2066 => (x"f8",x"87",x"ff",x"fd"),
  2067 => (x"26",x"87",x"c2",x"8e"),
  2068 => (x"26",x"4c",x"26",x"4d"),
  2069 => (x"0e",x"4f",x"26",x"4b"),
  2070 => (x"5d",x"5c",x"5b",x"5e"),
  2071 => (x"71",x"86",x"f8",x"0e"),
  2072 => (x"4c",x"a5",x"c4",x"4d"),
  2073 => (x"a8",x"6c",x"48",x"6d"),
  2074 => (x"ff",x"87",x"c5",x"05"),
  2075 => (x"87",x"e5",x"c0",x"48"),
  2076 => (x"d0",x"87",x"df",x"fd"),
  2077 => (x"48",x"6c",x"4b",x"a5"),
  2078 => (x"a6",x"c4",x"90",x"c4"),
  2079 => (x"6b",x"83",x"70",x"58"),
  2080 => (x"9b",x"ff",x"c3",x"4b"),
  2081 => (x"80",x"c1",x"48",x"6c"),
  2082 => (x"cf",x"58",x"a6",x"c8"),
  2083 => (x"fc",x"7c",x"70",x"98"),
  2084 => (x"49",x"73",x"87",x"f8"),
  2085 => (x"fe",x"8e",x"f8",x"48"),
  2086 => (x"73",x"1e",x"87",x"f5"),
  2087 => (x"fc",x"86",x"f8",x"1e"),
  2088 => (x"bf",x"e0",x"87",x"f0"),
  2089 => (x"e0",x"c0",x"49",x"4b"),
  2090 => (x"c0",x"02",x"99",x"c0"),
  2091 => (x"4a",x"73",x"87",x"e7"),
  2092 => (x"c3",x"9a",x"ff",x"c3"),
  2093 => (x"48",x"bf",x"fe",x"c1"),
  2094 => (x"a6",x"c4",x"90",x"c4"),
  2095 => (x"ce",x"c2",x"c3",x"58"),
  2096 => (x"72",x"81",x"70",x"49"),
  2097 => (x"fe",x"c1",x"c3",x"79"),
  2098 => (x"80",x"c1",x"48",x"bf"),
  2099 => (x"cf",x"58",x"a6",x"c8"),
  2100 => (x"c2",x"c2",x"c3",x"98"),
  2101 => (x"d0",x"49",x"73",x"58"),
  2102 => (x"c0",x"02",x"99",x"c0"),
  2103 => (x"c2",x"c3",x"87",x"f2"),
  2104 => (x"c3",x"48",x"bf",x"c6"),
  2105 => (x"a8",x"bf",x"ca",x"c2"),
  2106 => (x"87",x"e4",x"c0",x"02"),
  2107 => (x"bf",x"c6",x"c2",x"c3"),
  2108 => (x"c4",x"90",x"c4",x"48"),
  2109 => (x"c3",x"c3",x"58",x"a6"),
  2110 => (x"81",x"70",x"49",x"ce"),
  2111 => (x"78",x"69",x"48",x"e0"),
  2112 => (x"bf",x"c6",x"c2",x"c3"),
  2113 => (x"c8",x"80",x"c1",x"48"),
  2114 => (x"98",x"cf",x"58",x"a6"),
  2115 => (x"58",x"ca",x"c2",x"c3"),
  2116 => (x"c4",x"87",x"f0",x"fa"),
  2117 => (x"f1",x"fa",x"58",x"a6"),
  2118 => (x"fc",x"8e",x"f8",x"87"),
  2119 => (x"c3",x"1e",x"87",x"f5"),
  2120 => (x"fa",x"49",x"fe",x"c1"),
  2121 => (x"c2",x"c2",x"87",x"f4"),
  2122 => (x"c7",x"f9",x"49",x"da"),
  2123 => (x"87",x"f5",x"c3",x"87"),
  2124 => (x"73",x"1e",x"4f",x"26"),
  2125 => (x"fe",x"c1",x"c3",x"1e"),
  2126 => (x"87",x"db",x"fc",x"49"),
  2127 => (x"b7",x"c0",x"4a",x"70"),
  2128 => (x"cc",x"c2",x"04",x"aa"),
  2129 => (x"aa",x"f0",x"c3",x"87"),
  2130 => (x"c2",x"87",x"c9",x"05"),
  2131 => (x"c1",x"48",x"dd",x"c7"),
  2132 => (x"87",x"ed",x"c1",x"78"),
  2133 => (x"05",x"aa",x"e0",x"c3"),
  2134 => (x"c7",x"c2",x"87",x"c9"),
  2135 => (x"78",x"c1",x"48",x"e1"),
  2136 => (x"c2",x"87",x"de",x"c1"),
  2137 => (x"02",x"bf",x"e1",x"c7"),
  2138 => (x"c0",x"c2",x"87",x"c6"),
  2139 => (x"87",x"c2",x"4b",x"a2"),
  2140 => (x"c7",x"c2",x"4b",x"72"),
  2141 => (x"c0",x"02",x"bf",x"dd"),
  2142 => (x"49",x"73",x"87",x"e0"),
  2143 => (x"91",x"29",x"b7",x"c4"),
  2144 => (x"81",x"e5",x"c7",x"c2"),
  2145 => (x"9a",x"cf",x"4a",x"73"),
  2146 => (x"48",x"c1",x"92",x"c2"),
  2147 => (x"4a",x"70",x"30",x"72"),
  2148 => (x"48",x"72",x"ba",x"ff"),
  2149 => (x"79",x"70",x"98",x"69"),
  2150 => (x"49",x"73",x"87",x"db"),
  2151 => (x"91",x"29",x"b7",x"c4"),
  2152 => (x"81",x"e5",x"c7",x"c2"),
  2153 => (x"9a",x"cf",x"4a",x"73"),
  2154 => (x"48",x"c3",x"92",x"c2"),
  2155 => (x"4a",x"70",x"30",x"72"),
  2156 => (x"70",x"b0",x"69",x"48"),
  2157 => (x"e1",x"c7",x"c2",x"79"),
  2158 => (x"c2",x"78",x"c0",x"48"),
  2159 => (x"c0",x"48",x"dd",x"c7"),
  2160 => (x"fe",x"c1",x"c3",x"78"),
  2161 => (x"87",x"cf",x"fa",x"49"),
  2162 => (x"b7",x"c0",x"4a",x"70"),
  2163 => (x"f4",x"fd",x"03",x"aa"),
  2164 => (x"c4",x"48",x"c0",x"87"),
  2165 => (x"26",x"4d",x"26",x"87"),
  2166 => (x"26",x"4b",x"26",x"4c"),
  2167 => (x"00",x"00",x"00",x"4f"),
  2168 => (x"00",x"00",x"00",x"00"),
  2169 => (x"00",x"00",x"00",x"00"),
  2170 => (x"00",x"00",x"00",x"00"),
  2171 => (x"00",x"00",x"00",x"00"),
  2172 => (x"00",x"00",x"00",x"00"),
  2173 => (x"00",x"00",x"00",x"00"),
  2174 => (x"00",x"00",x"00",x"00"),
  2175 => (x"00",x"00",x"00",x"00"),
  2176 => (x"00",x"00",x"00",x"00"),
  2177 => (x"00",x"00",x"00",x"00"),
  2178 => (x"00",x"00",x"00",x"00"),
  2179 => (x"00",x"00",x"00",x"00"),
  2180 => (x"00",x"00",x"00",x"00"),
  2181 => (x"00",x"00",x"00",x"00"),
  2182 => (x"00",x"00",x"00",x"00"),
  2183 => (x"00",x"00",x"00",x"00"),
  2184 => (x"00",x"00",x"00",x"00"),
  2185 => (x"4a",x"c0",x"1e",x"00"),
  2186 => (x"91",x"c4",x"49",x"72"),
  2187 => (x"81",x"e5",x"c7",x"c2"),
  2188 => (x"82",x"c1",x"79",x"c0"),
  2189 => (x"04",x"aa",x"b7",x"d0"),
  2190 => (x"4f",x"26",x"87",x"ee"),
  2191 => (x"5c",x"5b",x"5e",x"0e"),
  2192 => (x"4d",x"71",x"0e",x"5d"),
  2193 => (x"75",x"87",x"cb",x"f6"),
  2194 => (x"2a",x"b7",x"c4",x"4a"),
  2195 => (x"e5",x"c7",x"c2",x"92"),
  2196 => (x"cf",x"4c",x"75",x"82"),
  2197 => (x"6a",x"94",x"c2",x"9c"),
  2198 => (x"2b",x"74",x"4b",x"49"),
  2199 => (x"48",x"c2",x"9b",x"c3"),
  2200 => (x"4c",x"70",x"30",x"74"),
  2201 => (x"48",x"74",x"bc",x"ff"),
  2202 => (x"7a",x"70",x"98",x"71"),
  2203 => (x"73",x"87",x"db",x"f5"),
  2204 => (x"87",x"e1",x"fd",x"48"),
  2205 => (x"d0",x"ff",x"1e",x"1e"),
  2206 => (x"c0",x"c8",x"48",x"bf"),
  2207 => (x"a6",x"c4",x"98",x"c0"),
  2208 => (x"02",x"98",x"70",x"58"),
  2209 => (x"d0",x"ff",x"87",x"d0"),
  2210 => (x"c0",x"c8",x"48",x"bf"),
  2211 => (x"a6",x"c4",x"98",x"c0"),
  2212 => (x"05",x"98",x"70",x"58"),
  2213 => (x"d0",x"ff",x"87",x"f0"),
  2214 => (x"78",x"e1",x"c4",x"48"),
  2215 => (x"d4",x"ff",x"48",x"71"),
  2216 => (x"66",x"c8",x"78",x"08"),
  2217 => (x"08",x"d4",x"ff",x"48"),
  2218 => (x"4f",x"26",x"26",x"78"),
  2219 => (x"4a",x"71",x"1e",x"1e"),
  2220 => (x"1e",x"49",x"66",x"c8"),
  2221 => (x"fb",x"fe",x"49",x"72"),
  2222 => (x"ff",x"86",x"c4",x"87"),
  2223 => (x"c8",x"48",x"bf",x"d0"),
  2224 => (x"c4",x"98",x"c0",x"c0"),
  2225 => (x"98",x"70",x"58",x"a6"),
  2226 => (x"ff",x"87",x"d0",x"02"),
  2227 => (x"c8",x"48",x"bf",x"d0"),
  2228 => (x"c4",x"98",x"c0",x"c0"),
  2229 => (x"98",x"70",x"58",x"a6"),
  2230 => (x"ff",x"87",x"f0",x"05"),
  2231 => (x"e0",x"c0",x"48",x"d0"),
  2232 => (x"4f",x"26",x"26",x"78"),
  2233 => (x"71",x"1e",x"73",x"1e"),
  2234 => (x"1e",x"66",x"c8",x"4b"),
  2235 => (x"e0",x"c1",x"4a",x"73"),
  2236 => (x"f7",x"fe",x"49",x"a2"),
  2237 => (x"87",x"c4",x"26",x"87"),
  2238 => (x"4c",x"26",x"4d",x"26"),
  2239 => (x"4f",x"26",x"4b",x"26"),
  2240 => (x"d0",x"ff",x"1e",x"1e"),
  2241 => (x"c0",x"c8",x"48",x"bf"),
  2242 => (x"a6",x"c4",x"98",x"c0"),
  2243 => (x"02",x"98",x"70",x"58"),
  2244 => (x"d0",x"ff",x"87",x"d0"),
  2245 => (x"c0",x"c8",x"48",x"bf"),
  2246 => (x"a6",x"c4",x"98",x"c0"),
  2247 => (x"05",x"98",x"70",x"58"),
  2248 => (x"d0",x"ff",x"87",x"f0"),
  2249 => (x"78",x"c9",x"c4",x"48"),
  2250 => (x"d4",x"ff",x"48",x"71"),
  2251 => (x"26",x"26",x"78",x"08"),
  2252 => (x"71",x"1e",x"1e",x"4f"),
  2253 => (x"c7",x"ff",x"49",x"4a"),
  2254 => (x"bf",x"d0",x"ff",x"87"),
  2255 => (x"c0",x"c0",x"c8",x"48"),
  2256 => (x"58",x"a6",x"c4",x"98"),
  2257 => (x"d0",x"02",x"98",x"70"),
  2258 => (x"bf",x"d0",x"ff",x"87"),
  2259 => (x"c0",x"c0",x"c8",x"48"),
  2260 => (x"58",x"a6",x"c4",x"98"),
  2261 => (x"f0",x"05",x"98",x"70"),
  2262 => (x"48",x"d0",x"ff",x"87"),
  2263 => (x"26",x"26",x"78",x"c8"),
  2264 => (x"1e",x"73",x"1e",x"4f"),
  2265 => (x"c3",x"4b",x"71",x"1e"),
  2266 => (x"02",x"bf",x"da",x"c4"),
  2267 => (x"cc",x"c3",x"87",x"c3"),
  2268 => (x"bf",x"d0",x"ff",x"87"),
  2269 => (x"c0",x"c0",x"c8",x"48"),
  2270 => (x"58",x"a6",x"c4",x"98"),
  2271 => (x"d0",x"02",x"98",x"70"),
  2272 => (x"bf",x"d0",x"ff",x"87"),
  2273 => (x"c0",x"c0",x"c8",x"48"),
  2274 => (x"58",x"a6",x"c4",x"98"),
  2275 => (x"f0",x"05",x"98",x"70"),
  2276 => (x"48",x"d0",x"ff",x"87"),
  2277 => (x"73",x"78",x"c9",x"c4"),
  2278 => (x"b0",x"e0",x"c0",x"48"),
  2279 => (x"78",x"08",x"d4",x"ff"),
  2280 => (x"48",x"ce",x"c4",x"c3"),
  2281 => (x"66",x"cc",x"78",x"c0"),
  2282 => (x"c3",x"87",x"c5",x"02"),
  2283 => (x"87",x"c2",x"49",x"ff"),
  2284 => (x"c4",x"c3",x"49",x"c0"),
  2285 => (x"66",x"d0",x"59",x"d6"),
  2286 => (x"c5",x"87",x"c6",x"02"),
  2287 => (x"c4",x"4a",x"d5",x"d5"),
  2288 => (x"ff",x"ff",x"cf",x"87"),
  2289 => (x"da",x"c4",x"c3",x"4a"),
  2290 => (x"da",x"c4",x"c3",x"5a"),
  2291 => (x"26",x"78",x"c1",x"48"),
  2292 => (x"4d",x"26",x"87",x"c4"),
  2293 => (x"4b",x"26",x"4c",x"26"),
  2294 => (x"5e",x"0e",x"4f",x"26"),
  2295 => (x"0e",x"5d",x"5c",x"5b"),
  2296 => (x"c4",x"c3",x"4a",x"71"),
  2297 => (x"72",x"4c",x"bf",x"d6"),
  2298 => (x"87",x"cb",x"02",x"9a"),
  2299 => (x"c2",x"91",x"c8",x"49"),
  2300 => (x"71",x"4b",x"db",x"ce"),
  2301 => (x"c2",x"87",x"c4",x"83"),
  2302 => (x"c0",x"4b",x"db",x"d2"),
  2303 => (x"74",x"49",x"13",x"4d"),
  2304 => (x"d2",x"c4",x"c3",x"99"),
  2305 => (x"b8",x"71",x"48",x"bf"),
  2306 => (x"78",x"08",x"d4",x"ff"),
  2307 => (x"85",x"2c",x"b7",x"c1"),
  2308 => (x"04",x"ad",x"b7",x"c8"),
  2309 => (x"c4",x"c3",x"87",x"e7"),
  2310 => (x"c8",x"48",x"bf",x"ce"),
  2311 => (x"d2",x"c4",x"c3",x"80"),
  2312 => (x"87",x"ee",x"fe",x"58"),
  2313 => (x"71",x"1e",x"73",x"1e"),
  2314 => (x"9a",x"4a",x"13",x"4b"),
  2315 => (x"72",x"87",x"cb",x"02"),
  2316 => (x"87",x"e6",x"fe",x"49"),
  2317 => (x"05",x"9a",x"4a",x"13"),
  2318 => (x"d9",x"fe",x"87",x"f5"),
  2319 => (x"c3",x"1e",x"1e",x"87"),
  2320 => (x"49",x"bf",x"ce",x"c4"),
  2321 => (x"48",x"ce",x"c4",x"c3"),
  2322 => (x"c4",x"78",x"a1",x"c1"),
  2323 => (x"03",x"a9",x"b7",x"c0"),
  2324 => (x"d4",x"ff",x"87",x"db"),
  2325 => (x"d2",x"c4",x"c3",x"48"),
  2326 => (x"c4",x"c3",x"78",x"bf"),
  2327 => (x"c3",x"49",x"bf",x"ce"),
  2328 => (x"c1",x"48",x"ce",x"c4"),
  2329 => (x"c0",x"c4",x"78",x"a1"),
  2330 => (x"e5",x"04",x"a9",x"b7"),
  2331 => (x"bf",x"d0",x"ff",x"87"),
  2332 => (x"c0",x"c0",x"c8",x"48"),
  2333 => (x"58",x"a6",x"c4",x"98"),
  2334 => (x"d0",x"02",x"98",x"70"),
  2335 => (x"bf",x"d0",x"ff",x"87"),
  2336 => (x"c0",x"c0",x"c8",x"48"),
  2337 => (x"58",x"a6",x"c4",x"98"),
  2338 => (x"f0",x"05",x"98",x"70"),
  2339 => (x"48",x"d0",x"ff",x"87"),
  2340 => (x"c4",x"c3",x"78",x"c8"),
  2341 => (x"78",x"c0",x"48",x"da"),
  2342 => (x"00",x"4f",x"26",x"26"),
  2343 => (x"00",x"00",x"00",x"00"),
  2344 => (x"00",x"00",x"00",x"00"),
  2345 => (x"5f",x"5f",x"00",x"00"),
  2346 => (x"00",x"00",x"00",x"00"),
  2347 => (x"03",x"00",x"03",x"03"),
  2348 => (x"14",x"00",x"00",x"03"),
  2349 => (x"7f",x"14",x"7f",x"7f"),
  2350 => (x"00",x"00",x"14",x"7f"),
  2351 => (x"6b",x"6b",x"2e",x"24"),
  2352 => (x"4c",x"00",x"12",x"3a"),
  2353 => (x"6c",x"18",x"36",x"6a"),
  2354 => (x"30",x"00",x"32",x"56"),
  2355 => (x"77",x"59",x"4f",x"7e"),
  2356 => (x"00",x"40",x"68",x"3a"),
  2357 => (x"03",x"07",x"04",x"00"),
  2358 => (x"00",x"00",x"00",x"00"),
  2359 => (x"63",x"3e",x"1c",x"00"),
  2360 => (x"00",x"00",x"00",x"41"),
  2361 => (x"3e",x"63",x"41",x"00"),
  2362 => (x"08",x"00",x"00",x"1c"),
  2363 => (x"1c",x"1c",x"3e",x"2a"),
  2364 => (x"00",x"08",x"2a",x"3e"),
  2365 => (x"3e",x"3e",x"08",x"08"),
  2366 => (x"00",x"00",x"08",x"08"),
  2367 => (x"60",x"e0",x"80",x"00"),
  2368 => (x"00",x"00",x"00",x"00"),
  2369 => (x"08",x"08",x"08",x"08"),
  2370 => (x"00",x"00",x"08",x"08"),
  2371 => (x"60",x"60",x"00",x"00"),
  2372 => (x"40",x"00",x"00",x"00"),
  2373 => (x"0c",x"18",x"30",x"60"),
  2374 => (x"00",x"01",x"03",x"06"),
  2375 => (x"4d",x"59",x"7f",x"3e"),
  2376 => (x"00",x"00",x"3e",x"7f"),
  2377 => (x"7f",x"7f",x"06",x"04"),
  2378 => (x"00",x"00",x"00",x"00"),
  2379 => (x"59",x"71",x"63",x"42"),
  2380 => (x"00",x"00",x"46",x"4f"),
  2381 => (x"49",x"49",x"63",x"22"),
  2382 => (x"18",x"00",x"36",x"7f"),
  2383 => (x"7f",x"13",x"16",x"1c"),
  2384 => (x"00",x"00",x"10",x"7f"),
  2385 => (x"45",x"45",x"67",x"27"),
  2386 => (x"00",x"00",x"39",x"7d"),
  2387 => (x"49",x"4b",x"7e",x"3c"),
  2388 => (x"00",x"00",x"30",x"79"),
  2389 => (x"79",x"71",x"01",x"01"),
  2390 => (x"00",x"00",x"07",x"0f"),
  2391 => (x"49",x"49",x"7f",x"36"),
  2392 => (x"00",x"00",x"36",x"7f"),
  2393 => (x"69",x"49",x"4f",x"06"),
  2394 => (x"00",x"00",x"1e",x"3f"),
  2395 => (x"66",x"66",x"00",x"00"),
  2396 => (x"00",x"00",x"00",x"00"),
  2397 => (x"66",x"e6",x"80",x"00"),
  2398 => (x"00",x"00",x"00",x"00"),
  2399 => (x"14",x"14",x"08",x"08"),
  2400 => (x"00",x"00",x"22",x"22"),
  2401 => (x"14",x"14",x"14",x"14"),
  2402 => (x"00",x"00",x"14",x"14"),
  2403 => (x"14",x"14",x"22",x"22"),
  2404 => (x"00",x"00",x"08",x"08"),
  2405 => (x"59",x"51",x"03",x"02"),
  2406 => (x"3e",x"00",x"06",x"0f"),
  2407 => (x"55",x"5d",x"41",x"7f"),
  2408 => (x"00",x"00",x"1e",x"1f"),
  2409 => (x"09",x"09",x"7f",x"7e"),
  2410 => (x"00",x"00",x"7e",x"7f"),
  2411 => (x"49",x"49",x"7f",x"7f"),
  2412 => (x"00",x"00",x"36",x"7f"),
  2413 => (x"41",x"63",x"3e",x"1c"),
  2414 => (x"00",x"00",x"41",x"41"),
  2415 => (x"63",x"41",x"7f",x"7f"),
  2416 => (x"00",x"00",x"1c",x"3e"),
  2417 => (x"49",x"49",x"7f",x"7f"),
  2418 => (x"00",x"00",x"41",x"41"),
  2419 => (x"09",x"09",x"7f",x"7f"),
  2420 => (x"00",x"00",x"01",x"01"),
  2421 => (x"49",x"41",x"7f",x"3e"),
  2422 => (x"00",x"00",x"7a",x"7b"),
  2423 => (x"08",x"08",x"7f",x"7f"),
  2424 => (x"00",x"00",x"7f",x"7f"),
  2425 => (x"7f",x"7f",x"41",x"00"),
  2426 => (x"00",x"00",x"00",x"41"),
  2427 => (x"40",x"40",x"60",x"20"),
  2428 => (x"7f",x"00",x"3f",x"7f"),
  2429 => (x"36",x"1c",x"08",x"7f"),
  2430 => (x"00",x"00",x"41",x"63"),
  2431 => (x"40",x"40",x"7f",x"7f"),
  2432 => (x"7f",x"00",x"40",x"40"),
  2433 => (x"06",x"0c",x"06",x"7f"),
  2434 => (x"7f",x"00",x"7f",x"7f"),
  2435 => (x"18",x"0c",x"06",x"7f"),
  2436 => (x"00",x"00",x"7f",x"7f"),
  2437 => (x"41",x"41",x"7f",x"3e"),
  2438 => (x"00",x"00",x"3e",x"7f"),
  2439 => (x"09",x"09",x"7f",x"7f"),
  2440 => (x"3e",x"00",x"06",x"0f"),
  2441 => (x"7f",x"61",x"41",x"7f"),
  2442 => (x"00",x"00",x"40",x"7e"),
  2443 => (x"19",x"09",x"7f",x"7f"),
  2444 => (x"00",x"00",x"66",x"7f"),
  2445 => (x"59",x"4d",x"6f",x"26"),
  2446 => (x"00",x"00",x"32",x"7b"),
  2447 => (x"7f",x"7f",x"01",x"01"),
  2448 => (x"00",x"00",x"01",x"01"),
  2449 => (x"40",x"40",x"7f",x"3f"),
  2450 => (x"00",x"00",x"3f",x"7f"),
  2451 => (x"70",x"70",x"3f",x"0f"),
  2452 => (x"7f",x"00",x"0f",x"3f"),
  2453 => (x"30",x"18",x"30",x"7f"),
  2454 => (x"41",x"00",x"7f",x"7f"),
  2455 => (x"1c",x"1c",x"36",x"63"),
  2456 => (x"01",x"41",x"63",x"36"),
  2457 => (x"7c",x"7c",x"06",x"03"),
  2458 => (x"61",x"01",x"03",x"06"),
  2459 => (x"47",x"4d",x"59",x"71"),
  2460 => (x"00",x"00",x"41",x"43"),
  2461 => (x"41",x"7f",x"7f",x"00"),
  2462 => (x"01",x"00",x"00",x"41"),
  2463 => (x"18",x"0c",x"06",x"03"),
  2464 => (x"00",x"40",x"60",x"30"),
  2465 => (x"7f",x"41",x"41",x"00"),
  2466 => (x"08",x"00",x"00",x"7f"),
  2467 => (x"06",x"03",x"06",x"0c"),
  2468 => (x"80",x"00",x"08",x"0c"),
  2469 => (x"80",x"80",x"80",x"80"),
  2470 => (x"00",x"00",x"80",x"80"),
  2471 => (x"07",x"03",x"00",x"00"),
  2472 => (x"00",x"00",x"00",x"04"),
  2473 => (x"54",x"54",x"74",x"20"),
  2474 => (x"00",x"00",x"78",x"7c"),
  2475 => (x"44",x"44",x"7f",x"7f"),
  2476 => (x"00",x"00",x"38",x"7c"),
  2477 => (x"44",x"44",x"7c",x"38"),
  2478 => (x"00",x"00",x"00",x"44"),
  2479 => (x"44",x"44",x"7c",x"38"),
  2480 => (x"00",x"00",x"7f",x"7f"),
  2481 => (x"54",x"54",x"7c",x"38"),
  2482 => (x"00",x"00",x"18",x"5c"),
  2483 => (x"05",x"7f",x"7e",x"04"),
  2484 => (x"00",x"00",x"00",x"05"),
  2485 => (x"a4",x"a4",x"bc",x"18"),
  2486 => (x"00",x"00",x"7c",x"fc"),
  2487 => (x"04",x"04",x"7f",x"7f"),
  2488 => (x"00",x"00",x"78",x"7c"),
  2489 => (x"7d",x"3d",x"00",x"00"),
  2490 => (x"00",x"00",x"00",x"40"),
  2491 => (x"fd",x"80",x"80",x"80"),
  2492 => (x"00",x"00",x"00",x"7d"),
  2493 => (x"38",x"10",x"7f",x"7f"),
  2494 => (x"00",x"00",x"44",x"6c"),
  2495 => (x"7f",x"3f",x"00",x"00"),
  2496 => (x"7c",x"00",x"00",x"40"),
  2497 => (x"0c",x"18",x"0c",x"7c"),
  2498 => (x"00",x"00",x"78",x"7c"),
  2499 => (x"04",x"04",x"7c",x"7c"),
  2500 => (x"00",x"00",x"78",x"7c"),
  2501 => (x"44",x"44",x"7c",x"38"),
  2502 => (x"00",x"00",x"38",x"7c"),
  2503 => (x"24",x"24",x"fc",x"fc"),
  2504 => (x"00",x"00",x"18",x"3c"),
  2505 => (x"24",x"24",x"3c",x"18"),
  2506 => (x"00",x"00",x"fc",x"fc"),
  2507 => (x"04",x"04",x"7c",x"7c"),
  2508 => (x"00",x"00",x"08",x"0c"),
  2509 => (x"54",x"54",x"5c",x"48"),
  2510 => (x"00",x"00",x"20",x"74"),
  2511 => (x"44",x"7f",x"3f",x"04"),
  2512 => (x"00",x"00",x"00",x"44"),
  2513 => (x"40",x"40",x"7c",x"3c"),
  2514 => (x"00",x"00",x"7c",x"7c"),
  2515 => (x"60",x"60",x"3c",x"1c"),
  2516 => (x"3c",x"00",x"1c",x"3c"),
  2517 => (x"60",x"30",x"60",x"7c"),
  2518 => (x"44",x"00",x"3c",x"7c"),
  2519 => (x"38",x"10",x"38",x"6c"),
  2520 => (x"00",x"00",x"44",x"6c"),
  2521 => (x"60",x"e0",x"bc",x"1c"),
  2522 => (x"00",x"00",x"1c",x"3c"),
  2523 => (x"5c",x"74",x"64",x"44"),
  2524 => (x"00",x"00",x"44",x"4c"),
  2525 => (x"77",x"3e",x"08",x"08"),
  2526 => (x"00",x"00",x"41",x"41"),
  2527 => (x"7f",x"7f",x"00",x"00"),
  2528 => (x"00",x"00",x"00",x"00"),
  2529 => (x"3e",x"77",x"41",x"41"),
  2530 => (x"02",x"00",x"08",x"08"),
  2531 => (x"02",x"03",x"01",x"01"),
  2532 => (x"7f",x"00",x"01",x"02"),
  2533 => (x"7f",x"7f",x"7f",x"7f"),
  2534 => (x"08",x"00",x"7f",x"7f"),
  2535 => (x"3e",x"1c",x"1c",x"08"),
  2536 => (x"7f",x"7f",x"7f",x"3e"),
  2537 => (x"1c",x"3e",x"3e",x"7f"),
  2538 => (x"00",x"08",x"08",x"1c"),
  2539 => (x"7c",x"7c",x"18",x"10"),
  2540 => (x"00",x"00",x"10",x"18"),
  2541 => (x"7c",x"7c",x"30",x"10"),
  2542 => (x"10",x"00",x"10",x"30"),
  2543 => (x"78",x"60",x"60",x"30"),
  2544 => (x"42",x"00",x"06",x"1e"),
  2545 => (x"3c",x"18",x"3c",x"66"),
  2546 => (x"78",x"00",x"42",x"66"),
  2547 => (x"c6",x"c2",x"6a",x"38"),
  2548 => (x"60",x"00",x"38",x"6c"),
  2549 => (x"00",x"60",x"00",x"00"),
  2550 => (x"0e",x"00",x"60",x"00"),
  2551 => (x"5d",x"5c",x"5b",x"5e"),
  2552 => (x"4c",x"71",x"1e",x"0e"),
  2553 => (x"bf",x"e2",x"c4",x"c3"),
  2554 => (x"e6",x"c4",x"c3",x"4b"),
  2555 => (x"74",x"78",x"c0",x"48"),
  2556 => (x"c6",x"e2",x"c2",x"1e"),
  2557 => (x"c3",x"e2",x"fd",x"1e"),
  2558 => (x"97",x"86",x"c8",x"87"),
  2559 => (x"02",x"99",x"49",x"6b"),
  2560 => (x"c0",x"87",x"c8",x"c1"),
  2561 => (x"e6",x"c4",x"c3",x"1e"),
  2562 => (x"ad",x"74",x"4d",x"bf"),
  2563 => (x"c4",x"87",x"c7",x"02"),
  2564 => (x"78",x"c0",x"48",x"a6"),
  2565 => (x"a6",x"c4",x"87",x"c5"),
  2566 => (x"c4",x"78",x"c1",x"48"),
  2567 => (x"49",x"75",x"1e",x"66"),
  2568 => (x"c8",x"87",x"fe",x"ec"),
  2569 => (x"49",x"e0",x"c0",x"86"),
  2570 => (x"c4",x"87",x"ef",x"ee"),
  2571 => (x"49",x"6a",x"4a",x"a3"),
  2572 => (x"f0",x"87",x"f1",x"ef"),
  2573 => (x"c4",x"c3",x"87",x"c7"),
  2574 => (x"c1",x"48",x"bf",x"e6"),
  2575 => (x"ea",x"c4",x"c3",x"80"),
  2576 => (x"97",x"83",x"cc",x"58"),
  2577 => (x"05",x"99",x"49",x"6b"),
  2578 => (x"c3",x"87",x"f8",x"fe"),
  2579 => (x"4d",x"bf",x"e6",x"c4"),
  2580 => (x"03",x"ad",x"b7",x"c8"),
  2581 => (x"1e",x"c0",x"87",x"d9"),
  2582 => (x"e6",x"c4",x"c3",x"1e"),
  2583 => (x"c0",x"ec",x"49",x"bf"),
  2584 => (x"ef",x"86",x"c8",x"87"),
  2585 => (x"85",x"c1",x"87",x"d7"),
  2586 => (x"04",x"ad",x"b7",x"c8"),
  2587 => (x"c3",x"87",x"e7",x"ff"),
  2588 => (x"1e",x"bf",x"e6",x"c4"),
  2589 => (x"1e",x"d8",x"e2",x"c2"),
  2590 => (x"87",x"c0",x"e0",x"fd"),
  2591 => (x"4d",x"26",x"8e",x"f4"),
  2592 => (x"4b",x"26",x"4c",x"26"),
  2593 => (x"69",x"48",x"4f",x"26"),
  2594 => (x"69",x"6c",x"68",x"67"),
  2595 => (x"20",x"74",x"68",x"67"),
  2596 => (x"20",x"77",x"6f",x"72"),
  2597 => (x"00",x"0a",x"64",x"25"),
  2598 => (x"75",x"6e",x"65",x"4d"),
  2599 => (x"73",x"61",x"68",x"20"),
  2600 => (x"20",x"64",x"25",x"20"),
  2601 => (x"73",x"77",x"6f",x"72"),
  2602 => (x"61",x"43",x"00",x"0a"),
  2603 => (x"61",x"62",x"6c",x"6c"),
  2604 => (x"25",x"20",x"6b",x"63"),
  2605 => (x"45",x"00",x"0a",x"78"),
  2606 => (x"72",x"65",x"74",x"6e"),
  2607 => (x"74",x"65",x"64",x"20"),
  2608 => (x"65",x"74",x"63",x"65"),
  2609 => (x"64",x"25",x"20",x"64"),
  2610 => (x"63",x"20",x"2d",x"20"),
  2611 => (x"65",x"72",x"72",x"75"),
  2612 => (x"6f",x"72",x"74",x"6e"),
  2613 => (x"64",x"25",x"20",x"77"),
  2614 => (x"71",x"1e",x"00",x"0a"),
  2615 => (x"e6",x"c4",x"c3",x"4a"),
  2616 => (x"ea",x"c4",x"c3",x"5a"),
  2617 => (x"f2",x"fb",x"49",x"bf"),
  2618 => (x"e6",x"c4",x"c3",x"87"),
  2619 => (x"89",x"c1",x"49",x"bf"),
  2620 => (x"59",x"ee",x"c4",x"c3"),
  2621 => (x"87",x"e3",x"fb",x"71"),
  2622 => (x"c1",x"1e",x"4f",x"26"),
  2623 => (x"f0",x"e8",x"49",x"c0"),
  2624 => (x"fc",x"ef",x"c2",x"87"),
  2625 => (x"26",x"78",x"c0",x"48"),
  2626 => (x"5b",x"5e",x"0e",x"4f"),
  2627 => (x"e8",x"0e",x"5d",x"5c"),
  2628 => (x"c0",x"c8",x"4c",x"bf"),
  2629 => (x"ef",x"c2",x"4d",x"c0"),
  2630 => (x"49",x"13",x"4b",x"e8"),
  2631 => (x"70",x"87",x"dd",x"e4"),
  2632 => (x"87",x"c2",x"02",x"98"),
  2633 => (x"b7",x"c1",x"b4",x"75"),
  2634 => (x"87",x"ee",x"05",x"2d"),
  2635 => (x"b7",x"c8",x"49",x"74"),
  2636 => (x"c0",x"1e",x"71",x"29"),
  2637 => (x"87",x"ec",x"e6",x"49"),
  2638 => (x"ff",x"c3",x"49",x"74"),
  2639 => (x"c1",x"1e",x"71",x"99"),
  2640 => (x"87",x"e0",x"e6",x"49"),
  2641 => (x"f5",x"fc",x"8e",x"f8"),
  2642 => (x"5b",x"5e",x"0e",x"87"),
  2643 => (x"f0",x"0e",x"5d",x"5c"),
  2644 => (x"48",x"a6",x"c8",x"86"),
  2645 => (x"80",x"c4",x"78",x"c0"),
  2646 => (x"bf",x"ec",x"78",x"c0"),
  2647 => (x"c3",x"80",x"f8",x"7e"),
  2648 => (x"78",x"bf",x"e2",x"c4"),
  2649 => (x"bf",x"ee",x"c4",x"c3"),
  2650 => (x"e3",x"49",x"c7",x"4c"),
  2651 => (x"49",x"70",x"87",x"ce"),
  2652 => (x"ce",x"05",x"99",x"c2"),
  2653 => (x"f8",x"ef",x"c2",x"87"),
  2654 => (x"b9",x"ff",x"49",x"bf"),
  2655 => (x"99",x"c1",x"99",x"6e"),
  2656 => (x"c2",x"87",x"d7",x"02"),
  2657 => (x"4a",x"bf",x"fc",x"ef"),
  2658 => (x"f0",x"c2",x"ba",x"c1"),
  2659 => (x"c0",x"c1",x"5a",x"c0"),
  2660 => (x"dc",x"e6",x"49",x"a2"),
  2661 => (x"48",x"a6",x"cc",x"87"),
  2662 => (x"ef",x"c2",x"78",x"c1"),
  2663 => (x"78",x"6e",x"48",x"f8"),
  2664 => (x"bf",x"fc",x"ef",x"c2"),
  2665 => (x"fd",x"87",x"d7",x"05"),
  2666 => (x"fd",x"c3",x"87",x"df"),
  2667 => (x"87",x"cc",x"e2",x"49"),
  2668 => (x"e2",x"49",x"fa",x"c3"),
  2669 => (x"ef",x"c2",x"87",x"c6"),
  2670 => (x"c8",x"48",x"bf",x"fc"),
  2671 => (x"f5",x"c3",x"87",x"e5"),
  2672 => (x"87",x"f8",x"e1",x"49"),
  2673 => (x"99",x"c2",x"49",x"70"),
  2674 => (x"87",x"ec",x"c0",x"02"),
  2675 => (x"bf",x"ea",x"c4",x"c3"),
  2676 => (x"48",x"87",x"c9",x"02"),
  2677 => (x"c4",x"c3",x"88",x"c1"),
  2678 => (x"87",x"d7",x"58",x"ee"),
  2679 => (x"bf",x"e6",x"c4",x"c3"),
  2680 => (x"c4",x"91",x"cc",x"49"),
  2681 => (x"a1",x"c8",x"81",x"66"),
  2682 => (x"02",x"bf",x"6e",x"7e"),
  2683 => (x"ff",x"4b",x"87",x"c5"),
  2684 => (x"cc",x"0f",x"73",x"49"),
  2685 => (x"78",x"c1",x"48",x"a6"),
  2686 => (x"e0",x"49",x"f2",x"c3"),
  2687 => (x"49",x"70",x"87",x"fe"),
  2688 => (x"c0",x"02",x"99",x"c2"),
  2689 => (x"a6",x"cc",x"87",x"fb"),
  2690 => (x"e6",x"c4",x"c3",x"48"),
  2691 => (x"66",x"cc",x"78",x"bf"),
  2692 => (x"c3",x"89",x"c1",x"49"),
  2693 => (x"7e",x"bf",x"ea",x"c4"),
  2694 => (x"06",x"a9",x"b7",x"6e"),
  2695 => (x"c1",x"48",x"87",x"c9"),
  2696 => (x"ee",x"c4",x"c3",x"80"),
  2697 => (x"cc",x"87",x"d5",x"58"),
  2698 => (x"91",x"cc",x"49",x"66"),
  2699 => (x"c8",x"81",x"66",x"c4"),
  2700 => (x"bf",x"6e",x"7e",x"a1"),
  2701 => (x"4b",x"87",x"c5",x"02"),
  2702 => (x"0f",x"73",x"49",x"fe"),
  2703 => (x"c1",x"48",x"a6",x"cc"),
  2704 => (x"49",x"fd",x"c3",x"78"),
  2705 => (x"87",x"f4",x"df",x"ff"),
  2706 => (x"99",x"c2",x"49",x"70"),
  2707 => (x"87",x"ed",x"c0",x"02"),
  2708 => (x"bf",x"ea",x"c4",x"c3"),
  2709 => (x"87",x"c8",x"c0",x"02"),
  2710 => (x"48",x"ea",x"c4",x"c3"),
  2711 => (x"87",x"d8",x"78",x"c0"),
  2712 => (x"bf",x"e6",x"c4",x"c3"),
  2713 => (x"c4",x"91",x"cc",x"49"),
  2714 => (x"a1",x"c8",x"81",x"66"),
  2715 => (x"02",x"bf",x"6e",x"7e"),
  2716 => (x"4b",x"87",x"c5",x"c0"),
  2717 => (x"0f",x"73",x"49",x"fd"),
  2718 => (x"c1",x"48",x"a6",x"cc"),
  2719 => (x"49",x"fa",x"c3",x"78"),
  2720 => (x"87",x"f8",x"de",x"ff"),
  2721 => (x"99",x"c2",x"49",x"70"),
  2722 => (x"87",x"ff",x"c0",x"02"),
  2723 => (x"c3",x"48",x"a6",x"cc"),
  2724 => (x"78",x"bf",x"e6",x"c4"),
  2725 => (x"c1",x"48",x"66",x"cc"),
  2726 => (x"58",x"a6",x"c4",x"88"),
  2727 => (x"bf",x"ea",x"c4",x"c3"),
  2728 => (x"a8",x"b7",x"6e",x"48"),
  2729 => (x"87",x"c8",x"c0",x"03"),
  2730 => (x"48",x"ea",x"c4",x"c3"),
  2731 => (x"87",x"d6",x"78",x"6e"),
  2732 => (x"cc",x"49",x"66",x"cc"),
  2733 => (x"81",x"66",x"c4",x"91"),
  2734 => (x"6e",x"7e",x"a1",x"c8"),
  2735 => (x"c5",x"c0",x"02",x"bf"),
  2736 => (x"49",x"fc",x"4b",x"87"),
  2737 => (x"a6",x"cc",x"0f",x"73"),
  2738 => (x"c3",x"78",x"c1",x"48"),
  2739 => (x"4b",x"bf",x"ea",x"c4"),
  2740 => (x"06",x"ab",x"b7",x"c0"),
  2741 => (x"c1",x"87",x"c9",x"c0"),
  2742 => (x"ab",x"b7",x"c0",x"8b"),
  2743 => (x"87",x"f7",x"ff",x"01"),
  2744 => (x"ff",x"49",x"da",x"c1"),
  2745 => (x"70",x"87",x"d5",x"dd"),
  2746 => (x"9b",x"c2",x"4b",x"49"),
  2747 => (x"c2",x"02",x"9b",x"73"),
  2748 => (x"c4",x"c3",x"87",x"f1"),
  2749 => (x"c3",x"4d",x"bf",x"e2"),
  2750 => (x"1e",x"bf",x"ea",x"c4"),
  2751 => (x"e2",x"c2",x"1e",x"73"),
  2752 => (x"d5",x"fd",x"1e",x"f7"),
  2753 => (x"86",x"cc",x"87",x"f6"),
  2754 => (x"bf",x"ea",x"c4",x"c3"),
  2755 => (x"ab",x"b7",x"c0",x"4b"),
  2756 => (x"87",x"cb",x"c0",x"06"),
  2757 => (x"8b",x"c1",x"85",x"cc"),
  2758 => (x"01",x"ab",x"b7",x"c0"),
  2759 => (x"97",x"87",x"f5",x"ff"),
  2760 => (x"8a",x"c1",x"4a",x"6d"),
  2761 => (x"87",x"f5",x"c0",x"02"),
  2762 => (x"d5",x"c0",x"02",x"8a"),
  2763 => (x"c1",x"02",x"8a",x"87"),
  2764 => (x"05",x"8a",x"87",x"cb"),
  2765 => (x"c8",x"87",x"ec",x"c1"),
  2766 => (x"49",x"6a",x"4a",x"a5"),
  2767 => (x"c1",x"87",x"db",x"f6"),
  2768 => (x"a5",x"c8",x"87",x"e1"),
  2769 => (x"c2",x"1e",x"6b",x"4b"),
  2770 => (x"fd",x"1e",x"ea",x"e2"),
  2771 => (x"c8",x"87",x"ed",x"d4"),
  2772 => (x"c3",x"4b",x"6b",x"86"),
  2773 => (x"49",x"bf",x"ea",x"c4"),
  2774 => (x"c6",x"c1",x"0f",x"73"),
  2775 => (x"49",x"a5",x"c8",x"87"),
  2776 => (x"30",x"69",x"48",x"c1"),
  2777 => (x"c4",x"c3",x"49",x"70"),
  2778 => (x"71",x"48",x"bf",x"de"),
  2779 => (x"e2",x"c4",x"c3",x"b8"),
  2780 => (x"48",x"a6",x"cc",x"58"),
  2781 => (x"80",x"fc",x"78",x"c1"),
  2782 => (x"e6",x"c0",x"78",x"c1"),
  2783 => (x"49",x"a5",x"c8",x"87"),
  2784 => (x"6e",x"7e",x"a5",x"cb"),
  2785 => (x"c1",x"4a",x"bf",x"97"),
  2786 => (x"69",x"97",x"4b",x"a2"),
  2787 => (x"04",x"ab",x"b7",x"49"),
  2788 => (x"c0",x"87",x"c2",x"c0"),
  2789 => (x"97",x"0b",x"6e",x"4b"),
  2790 => (x"a6",x"cc",x"0b",x"7b"),
  2791 => (x"fc",x"78",x"c1",x"48"),
  2792 => (x"74",x"78",x"c1",x"80"),
  2793 => (x"e9",x"c0",x"02",x"9c"),
  2794 => (x"c0",x"02",x"6c",x"87"),
  2795 => (x"49",x"6c",x"87",x"e4"),
  2796 => (x"87",x"c8",x"da",x"ff"),
  2797 => (x"99",x"c1",x"49",x"70"),
  2798 => (x"87",x"cb",x"c0",x"02"),
  2799 => (x"c3",x"4b",x"a4",x"c4"),
  2800 => (x"49",x"bf",x"ea",x"c4"),
  2801 => (x"c8",x"0f",x"4b",x"6b"),
  2802 => (x"c5",x"c0",x"02",x"84"),
  2803 => (x"ff",x"05",x"6c",x"87"),
  2804 => (x"66",x"cc",x"87",x"dc"),
  2805 => (x"87",x"c8",x"c0",x"02"),
  2806 => (x"bf",x"ea",x"c4",x"c3"),
  2807 => (x"87",x"fb",x"ef",x"49"),
  2808 => (x"f0",x"48",x"66",x"c8"),
  2809 => (x"87",x"d6",x"f2",x"8e"),
  2810 => (x"14",x"91",x"12",x"58"),
  2811 => (x"23",x"1c",x"1b",x"1d"),
  2812 => (x"91",x"94",x"59",x"5a"),
  2813 => (x"f4",x"eb",x"f2",x"f5"),
  2814 => (x"00",x"00",x"00",x"00"),
  2815 => (x"00",x"00",x"00",x"00"),
  2816 => (x"00",x"00",x"1f",x"b1"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

