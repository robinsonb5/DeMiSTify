
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"c1",x"c3",x"87"),
    12 => (x"86",x"c0",x"d0",x"4e"),
    13 => (x"49",x"c0",x"c1",x"c3"),
    14 => (x"48",x"cc",x"ec",x"c2"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"cc",x"ec",x"c2",x"87"),
    21 => (x"c8",x"ec",x"c2",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"f3",x"c1",x"87",x"f7"),
    25 => (x"ec",x"c2",x"87",x"d5"),
    26 => (x"ec",x"c2",x"4d",x"cc"),
    27 => (x"ad",x"74",x"4c",x"cc"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"5c",x"5b",x"5e",x"0e"),
    32 => (x"86",x"f0",x"0e",x"5d"),
    33 => (x"a6",x"c4",x"4c",x"c0"),
    34 => (x"c0",x"78",x"c0",x"48"),
    35 => (x"c0",x"4b",x"a6",x"e4"),
    36 => (x"48",x"49",x"66",x"e0"),
    37 => (x"e4",x"c0",x"80",x"c1"),
    38 => (x"48",x"11",x"58",x"a6"),
    39 => (x"70",x"58",x"a6",x"c4"),
    40 => (x"f6",x"c3",x"02",x"98"),
    41 => (x"02",x"66",x"c4",x"87"),
    42 => (x"c4",x"87",x"c6",x"c3"),
    43 => (x"78",x"c0",x"48",x"a6"),
    44 => (x"f0",x"c0",x"4a",x"6e"),
    45 => (x"da",x"c2",x"02",x"8a"),
    46 => (x"8a",x"f3",x"c0",x"87"),
    47 => (x"87",x"db",x"c2",x"02"),
    48 => (x"dc",x"02",x"8a",x"c1"),
    49 => (x"02",x"8a",x"c8",x"87"),
    50 => (x"c4",x"87",x"c8",x"c2"),
    51 => (x"87",x"d1",x"02",x"8a"),
    52 => (x"c1",x"02",x"8a",x"c3"),
    53 => (x"8a",x"c2",x"87",x"eb"),
    54 => (x"c3",x"87",x"c6",x"02"),
    55 => (x"c9",x"c2",x"05",x"8a"),
    56 => (x"73",x"83",x"c4",x"87"),
    57 => (x"69",x"89",x"c4",x"49"),
    58 => (x"c1",x"02",x"6e",x"7e"),
    59 => (x"a6",x"c8",x"87",x"c8"),
    60 => (x"c4",x"78",x"c0",x"48"),
    61 => (x"cc",x"78",x"c0",x"80"),
    62 => (x"4a",x"6e",x"4d",x"66"),
    63 => (x"cf",x"2a",x"b7",x"dc"),
    64 => (x"c4",x"48",x"6e",x"9a"),
    65 => (x"72",x"58",x"a6",x"30"),
    66 => (x"87",x"c5",x"02",x"9a"),
    67 => (x"c1",x"48",x"a6",x"c8"),
    68 => (x"06",x"aa",x"c9",x"78"),
    69 => (x"f7",x"c0",x"87",x"c5"),
    70 => (x"c0",x"87",x"c3",x"82"),
    71 => (x"66",x"c8",x"82",x"f0"),
    72 => (x"72",x"87",x"c7",x"02"),
    73 => (x"87",x"f3",x"c2",x"49"),
    74 => (x"85",x"c1",x"84",x"c1"),
    75 => (x"04",x"ad",x"b7",x"c8"),
    76 => (x"c1",x"87",x"c7",x"ff"),
    77 => (x"f0",x"c0",x"87",x"cf"),
    78 => (x"87",x"df",x"c2",x"49"),
    79 => (x"c4",x"c1",x"84",x"c1"),
    80 => (x"73",x"83",x"c4",x"87"),
    81 => (x"6a",x"8a",x"c4",x"4a"),
    82 => (x"87",x"db",x"c1",x"49"),
    83 => (x"4c",x"a4",x"49",x"70"),
    84 => (x"c4",x"87",x"f2",x"c0"),
    85 => (x"78",x"c1",x"48",x"a6"),
    86 => (x"c4",x"87",x"ea",x"c0"),
    87 => (x"c4",x"4a",x"73",x"83"),
    88 => (x"c1",x"49",x"6a",x"8a"),
    89 => (x"84",x"c1",x"87",x"f5"),
    90 => (x"49",x"6e",x"87",x"db"),
    91 => (x"d4",x"87",x"ec",x"c1"),
    92 => (x"c0",x"48",x"6e",x"87"),
    93 => (x"c7",x"05",x"a8",x"e5"),
    94 => (x"48",x"a6",x"c4",x"87"),
    95 => (x"87",x"c5",x"78",x"c1"),
    96 => (x"d6",x"c1",x"49",x"6e"),
    97 => (x"66",x"e0",x"c0",x"87"),
    98 => (x"80",x"c1",x"48",x"49"),
    99 => (x"58",x"a6",x"e4",x"c0"),
   100 => (x"a6",x"c4",x"48",x"11"),
   101 => (x"05",x"98",x"70",x"58"),
   102 => (x"74",x"87",x"ca",x"fc"),
   103 => (x"26",x"8e",x"f0",x"48"),
   104 => (x"26",x"4c",x"26",x"4d"),
   105 => (x"0e",x"4f",x"26",x"4b"),
   106 => (x"0e",x"5c",x"5b",x"5e"),
   107 => (x"4c",x"c0",x"4b",x"71"),
   108 => (x"02",x"9a",x"4a",x"13"),
   109 => (x"49",x"72",x"87",x"cd"),
   110 => (x"c1",x"87",x"e0",x"c0"),
   111 => (x"9a",x"4a",x"13",x"84"),
   112 => (x"74",x"87",x"f3",x"05"),
   113 => (x"26",x"4c",x"26",x"48"),
   114 => (x"1e",x"4f",x"26",x"4b"),
   115 => (x"73",x"81",x"48",x"73"),
   116 => (x"87",x"c5",x"02",x"a9"),
   117 => (x"f6",x"05",x"53",x"12"),
   118 => (x"1e",x"4f",x"26",x"87"),
   119 => (x"4a",x"c0",x"ff",x"1e"),
   120 => (x"c0",x"c4",x"48",x"6a"),
   121 => (x"58",x"a6",x"c4",x"98"),
   122 => (x"f3",x"02",x"98",x"70"),
   123 => (x"48",x"7a",x"71",x"87"),
   124 => (x"1e",x"4f",x"26",x"26"),
   125 => (x"d4",x"ff",x"1e",x"73"),
   126 => (x"7b",x"ff",x"c3",x"4b"),
   127 => (x"ff",x"c3",x"4a",x"6b"),
   128 => (x"c8",x"49",x"6b",x"7b"),
   129 => (x"c3",x"b1",x"72",x"32"),
   130 => (x"4a",x"6b",x"7b",x"ff"),
   131 => (x"b2",x"71",x"31",x"c8"),
   132 => (x"6b",x"7b",x"ff",x"c3"),
   133 => (x"72",x"32",x"c8",x"49"),
   134 => (x"c4",x"48",x"71",x"b1"),
   135 => (x"26",x"4d",x"26",x"87"),
   136 => (x"26",x"4b",x"26",x"4c"),
   137 => (x"5b",x"5e",x"0e",x"4f"),
   138 => (x"71",x"0e",x"5d",x"5c"),
   139 => (x"4c",x"d4",x"ff",x"4a"),
   140 => (x"ff",x"c3",x"48",x"72"),
   141 => (x"c2",x"7c",x"70",x"98"),
   142 => (x"05",x"bf",x"cc",x"ec"),
   143 => (x"66",x"d0",x"87",x"c8"),
   144 => (x"d4",x"30",x"c9",x"48"),
   145 => (x"66",x"d0",x"58",x"a6"),
   146 => (x"71",x"29",x"d8",x"49"),
   147 => (x"98",x"ff",x"c3",x"48"),
   148 => (x"66",x"d0",x"7c",x"70"),
   149 => (x"71",x"29",x"d0",x"49"),
   150 => (x"98",x"ff",x"c3",x"48"),
   151 => (x"66",x"d0",x"7c",x"70"),
   152 => (x"71",x"29",x"c8",x"49"),
   153 => (x"98",x"ff",x"c3",x"48"),
   154 => (x"66",x"d0",x"7c",x"70"),
   155 => (x"98",x"ff",x"c3",x"48"),
   156 => (x"49",x"72",x"7c",x"70"),
   157 => (x"48",x"71",x"29",x"d0"),
   158 => (x"70",x"98",x"ff",x"c3"),
   159 => (x"c9",x"4b",x"6c",x"7c"),
   160 => (x"c3",x"4d",x"ff",x"f0"),
   161 => (x"d0",x"05",x"ab",x"ff"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"8d",x"c1",x"4b",x"6c"),
   164 => (x"c3",x"87",x"c6",x"02"),
   165 => (x"f0",x"02",x"ab",x"ff"),
   166 => (x"fd",x"48",x"73",x"87"),
   167 => (x"c0",x"1e",x"87",x"ff"),
   168 => (x"48",x"d4",x"ff",x"49"),
   169 => (x"c1",x"78",x"ff",x"c3"),
   170 => (x"b7",x"c8",x"c3",x"81"),
   171 => (x"87",x"f1",x"04",x"a9"),
   172 => (x"73",x"1e",x"4f",x"26"),
   173 => (x"c4",x"87",x"e7",x"1e"),
   174 => (x"c0",x"4b",x"df",x"f8"),
   175 => (x"f0",x"ff",x"c0",x"1e"),
   176 => (x"fd",x"49",x"f7",x"c1"),
   177 => (x"86",x"c4",x"87",x"df"),
   178 => (x"c0",x"05",x"a8",x"c1"),
   179 => (x"d4",x"ff",x"87",x"ea"),
   180 => (x"78",x"ff",x"c3",x"48"),
   181 => (x"c0",x"c0",x"c0",x"c1"),
   182 => (x"c0",x"1e",x"c0",x"c0"),
   183 => (x"e9",x"c1",x"f0",x"e1"),
   184 => (x"87",x"c1",x"fd",x"49"),
   185 => (x"98",x"70",x"86",x"c4"),
   186 => (x"ff",x"87",x"ca",x"05"),
   187 => (x"ff",x"c3",x"48",x"d4"),
   188 => (x"cb",x"48",x"c1",x"78"),
   189 => (x"87",x"e6",x"fe",x"87"),
   190 => (x"fe",x"05",x"8b",x"c1"),
   191 => (x"48",x"c0",x"87",x"fd"),
   192 => (x"1e",x"87",x"de",x"fc"),
   193 => (x"d4",x"ff",x"1e",x"73"),
   194 => (x"78",x"ff",x"c3",x"48"),
   195 => (x"fa",x"49",x"fe",x"cc"),
   196 => (x"4b",x"d3",x"87",x"d5"),
   197 => (x"ff",x"c0",x"1e",x"c0"),
   198 => (x"49",x"c1",x"c1",x"f0"),
   199 => (x"c4",x"87",x"c6",x"fc"),
   200 => (x"05",x"98",x"70",x"86"),
   201 => (x"d4",x"ff",x"87",x"ca"),
   202 => (x"78",x"ff",x"c3",x"48"),
   203 => (x"87",x"cb",x"48",x"c1"),
   204 => (x"c1",x"87",x"eb",x"fd"),
   205 => (x"db",x"ff",x"05",x"8b"),
   206 => (x"fb",x"48",x"c0",x"87"),
   207 => (x"4d",x"43",x"87",x"e3"),
   208 => (x"4d",x"43",x"00",x"44"),
   209 => (x"20",x"38",x"35",x"44"),
   210 => (x"20",x"0a",x"64",x"25"),
   211 => (x"4d",x"43",x"00",x"20"),
   212 => (x"5f",x"38",x"35",x"44"),
   213 => (x"64",x"25",x"20",x"32"),
   214 => (x"00",x"20",x"20",x"0a"),
   215 => (x"35",x"44",x"4d",x"43"),
   216 => (x"64",x"25",x"20",x"38"),
   217 => (x"00",x"20",x"20",x"0a"),
   218 => (x"43",x"48",x"44",x"53"),
   219 => (x"69",x"6e",x"49",x"20"),
   220 => (x"6c",x"61",x"69",x"74"),
   221 => (x"74",x"61",x"7a",x"69"),
   222 => (x"20",x"6e",x"6f",x"69"),
   223 => (x"6f",x"72",x"72",x"65"),
   224 => (x"00",x"0a",x"21",x"72"),
   225 => (x"5f",x"64",x"6d",x"63"),
   226 => (x"38",x"44",x"4d",x"43"),
   227 => (x"73",x"65",x"72",x"20"),
   228 => (x"73",x"6e",x"6f",x"70"),
   229 => (x"25",x"20",x"3a",x"65"),
   230 => (x"49",x"00",x"0a",x"64"),
   231 => (x"00",x"52",x"52",x"45"),
   232 => (x"00",x"49",x"50",x"53"),
   233 => (x"63",x"20",x"44",x"53"),
   234 => (x"20",x"64",x"72",x"61"),
   235 => (x"65",x"7a",x"69",x"73"),
   236 => (x"20",x"73",x"69",x"20"),
   237 => (x"00",x"0a",x"64",x"25"),
   238 => (x"74",x"69",x"72",x"57"),
   239 => (x"61",x"66",x"20",x"65"),
   240 => (x"64",x"65",x"6c",x"69"),
   241 => (x"5f",x"63",x"00",x"0a"),
   242 => (x"65",x"7a",x"69",x"73"),
   243 => (x"6c",x"75",x"6d",x"5f"),
   244 => (x"25",x"20",x"3a",x"74"),
   245 => (x"72",x"20",x"2c",x"64"),
   246 => (x"5f",x"64",x"61",x"65"),
   247 => (x"6c",x"5f",x"6c",x"62"),
   248 => (x"20",x"3a",x"6e",x"65"),
   249 => (x"20",x"2c",x"64",x"25"),
   250 => (x"7a",x"69",x"73",x"63"),
   251 => (x"25",x"20",x"3a",x"65"),
   252 => (x"4d",x"00",x"0a",x"64"),
   253 => (x"20",x"74",x"6c",x"75"),
   254 => (x"00",x"0a",x"64",x"25"),
   255 => (x"62",x"20",x"64",x"25"),
   256 => (x"6b",x"63",x"6f",x"6c"),
   257 => (x"66",x"6f",x"20",x"73"),
   258 => (x"7a",x"69",x"73",x"20"),
   259 => (x"64",x"25",x"20",x"65"),
   260 => (x"64",x"25",x"00",x"0a"),
   261 => (x"6f",x"6c",x"62",x"20"),
   262 => (x"20",x"73",x"6b",x"63"),
   263 => (x"35",x"20",x"66",x"6f"),
   264 => (x"62",x"20",x"32",x"31"),
   265 => (x"73",x"65",x"74",x"79"),
   266 => (x"5e",x"0e",x"00",x"0a"),
   267 => (x"0e",x"5d",x"5c",x"5b"),
   268 => (x"f9",x"4d",x"d4",x"ff"),
   269 => (x"ea",x"c6",x"87",x"e8"),
   270 => (x"f0",x"e1",x"c0",x"1e"),
   271 => (x"f7",x"49",x"c8",x"c1"),
   272 => (x"4b",x"70",x"87",x"e3"),
   273 => (x"1e",x"c4",x"ce",x"1e"),
   274 => (x"cc",x"87",x"f1",x"f0"),
   275 => (x"02",x"ab",x"c1",x"86"),
   276 => (x"ee",x"fa",x"87",x"c8"),
   277 => (x"c2",x"48",x"c0",x"87"),
   278 => (x"d6",x"f6",x"87",x"ca"),
   279 => (x"cf",x"49",x"70",x"87"),
   280 => (x"c6",x"99",x"ff",x"ff"),
   281 => (x"c8",x"02",x"a9",x"ea"),
   282 => (x"87",x"d7",x"fa",x"87"),
   283 => (x"f3",x"c1",x"48",x"c0"),
   284 => (x"7d",x"ff",x"c3",x"87"),
   285 => (x"f8",x"4c",x"f1",x"c0"),
   286 => (x"98",x"70",x"87",x"f8"),
   287 => (x"87",x"cb",x"c1",x"02"),
   288 => (x"ff",x"c0",x"1e",x"c0"),
   289 => (x"49",x"fa",x"c1",x"f0"),
   290 => (x"c4",x"87",x"da",x"f6"),
   291 => (x"9b",x"4b",x"70",x"86"),
   292 => (x"87",x"ed",x"c0",x"05"),
   293 => (x"1e",x"c2",x"cd",x"1e"),
   294 => (x"c3",x"87",x"e1",x"ef"),
   295 => (x"4b",x"6d",x"7d",x"ff"),
   296 => (x"1e",x"ce",x"cd",x"1e"),
   297 => (x"d0",x"87",x"d5",x"ef"),
   298 => (x"7d",x"ff",x"c3",x"86"),
   299 => (x"73",x"7d",x"7d",x"7d"),
   300 => (x"99",x"c0",x"c1",x"49"),
   301 => (x"c1",x"87",x"c5",x"02"),
   302 => (x"87",x"e8",x"c0",x"48"),
   303 => (x"e3",x"c0",x"48",x"c0"),
   304 => (x"cd",x"1e",x"73",x"87"),
   305 => (x"f3",x"ee",x"1e",x"dc"),
   306 => (x"c2",x"86",x"c8",x"87"),
   307 => (x"87",x"cc",x"05",x"ac"),
   308 => (x"ee",x"1e",x"e8",x"cd"),
   309 => (x"86",x"c4",x"87",x"e6"),
   310 => (x"87",x"c8",x"48",x"c0"),
   311 => (x"fe",x"05",x"8c",x"c1"),
   312 => (x"48",x"c0",x"87",x"d5"),
   313 => (x"0e",x"87",x"f6",x"f4"),
   314 => (x"5d",x"5c",x"5b",x"5e"),
   315 => (x"d0",x"ff",x"1e",x"0e"),
   316 => (x"c0",x"c0",x"c8",x"4d"),
   317 => (x"cc",x"ec",x"c2",x"4b"),
   318 => (x"ce",x"78",x"c1",x"48"),
   319 => (x"e6",x"f2",x"49",x"e0"),
   320 => (x"6d",x"4c",x"c7",x"87"),
   321 => (x"c4",x"98",x"73",x"48"),
   322 => (x"98",x"70",x"58",x"a6"),
   323 => (x"6d",x"87",x"cc",x"02"),
   324 => (x"c4",x"98",x"73",x"48"),
   325 => (x"98",x"70",x"58",x"a6"),
   326 => (x"c2",x"87",x"f4",x"05"),
   327 => (x"87",x"fe",x"f5",x"7d"),
   328 => (x"98",x"73",x"48",x"6d"),
   329 => (x"70",x"58",x"a6",x"c4"),
   330 => (x"87",x"cc",x"02",x"98"),
   331 => (x"98",x"73",x"48",x"6d"),
   332 => (x"70",x"58",x"a6",x"c4"),
   333 => (x"87",x"f4",x"05",x"98"),
   334 => (x"1e",x"c0",x"7d",x"c3"),
   335 => (x"c1",x"d0",x"e5",x"c0"),
   336 => (x"e0",x"f3",x"49",x"c0"),
   337 => (x"c1",x"86",x"c4",x"87"),
   338 => (x"87",x"c1",x"05",x"a8"),
   339 => (x"05",x"ac",x"c2",x"4c"),
   340 => (x"db",x"ce",x"87",x"cb"),
   341 => (x"87",x"cf",x"f1",x"49"),
   342 => (x"d8",x"c1",x"48",x"c0"),
   343 => (x"05",x"8c",x"c1",x"87"),
   344 => (x"fb",x"87",x"e0",x"fe"),
   345 => (x"ec",x"c2",x"87",x"c4"),
   346 => (x"98",x"70",x"58",x"d0"),
   347 => (x"c1",x"87",x"cd",x"05"),
   348 => (x"f0",x"ff",x"c0",x"1e"),
   349 => (x"f2",x"49",x"d0",x"c1"),
   350 => (x"86",x"c4",x"87",x"eb"),
   351 => (x"c3",x"48",x"d4",x"ff"),
   352 => (x"e7",x"c5",x"78",x"ff"),
   353 => (x"d4",x"ec",x"c2",x"87"),
   354 => (x"ce",x"1e",x"70",x"58"),
   355 => (x"eb",x"eb",x"1e",x"e4"),
   356 => (x"6d",x"86",x"c8",x"87"),
   357 => (x"c4",x"98",x"73",x"48"),
   358 => (x"98",x"70",x"58",x"a6"),
   359 => (x"6d",x"87",x"cc",x"02"),
   360 => (x"c4",x"98",x"73",x"48"),
   361 => (x"98",x"70",x"58",x"a6"),
   362 => (x"c2",x"87",x"f4",x"05"),
   363 => (x"48",x"d4",x"ff",x"7d"),
   364 => (x"c1",x"78",x"ff",x"c3"),
   365 => (x"e4",x"f1",x"26",x"48"),
   366 => (x"5b",x"5e",x"0e",x"87"),
   367 => (x"1e",x"0e",x"5d",x"5c"),
   368 => (x"4b",x"c0",x"c0",x"c8"),
   369 => (x"ee",x"c5",x"4c",x"c0"),
   370 => (x"c4",x"4a",x"df",x"cd"),
   371 => (x"d4",x"ff",x"5c",x"a6"),
   372 => (x"7c",x"ff",x"c3",x"4c"),
   373 => (x"fe",x"c3",x"48",x"6c"),
   374 => (x"c0",x"c2",x"05",x"a8"),
   375 => (x"05",x"99",x"71",x"87"),
   376 => (x"ff",x"87",x"e2",x"c0"),
   377 => (x"73",x"48",x"bf",x"d0"),
   378 => (x"58",x"a6",x"c4",x"98"),
   379 => (x"ce",x"02",x"98",x"70"),
   380 => (x"bf",x"d0",x"ff",x"87"),
   381 => (x"c4",x"98",x"73",x"48"),
   382 => (x"98",x"70",x"58",x"a6"),
   383 => (x"ff",x"87",x"f2",x"05"),
   384 => (x"d1",x"c4",x"48",x"d0"),
   385 => (x"48",x"66",x"d4",x"78"),
   386 => (x"06",x"a8",x"b7",x"c0"),
   387 => (x"c3",x"87",x"e0",x"c0"),
   388 => (x"4a",x"6c",x"7c",x"ff"),
   389 => (x"c7",x"02",x"99",x"71"),
   390 => (x"97",x"0a",x"71",x"87"),
   391 => (x"81",x"c1",x"0a",x"7a"),
   392 => (x"c1",x"48",x"66",x"d4"),
   393 => (x"58",x"a6",x"d8",x"88"),
   394 => (x"01",x"a8",x"b7",x"c0"),
   395 => (x"c3",x"87",x"e0",x"ff"),
   396 => (x"71",x"7c",x"7c",x"ff"),
   397 => (x"e1",x"c0",x"05",x"99"),
   398 => (x"bf",x"d0",x"ff",x"87"),
   399 => (x"c4",x"98",x"73",x"48"),
   400 => (x"98",x"70",x"58",x"a6"),
   401 => (x"ff",x"87",x"ce",x"02"),
   402 => (x"73",x"48",x"bf",x"d0"),
   403 => (x"58",x"a6",x"c4",x"98"),
   404 => (x"f2",x"05",x"98",x"70"),
   405 => (x"48",x"d0",x"ff",x"87"),
   406 => (x"4a",x"c1",x"78",x"d0"),
   407 => (x"05",x"8a",x"c1",x"7e"),
   408 => (x"6e",x"87",x"ee",x"fd"),
   409 => (x"f4",x"ee",x"26",x"48"),
   410 => (x"5b",x"5e",x"0e",x"87"),
   411 => (x"71",x"1e",x"0e",x"5c"),
   412 => (x"c0",x"c0",x"c8",x"4a"),
   413 => (x"ff",x"4c",x"c0",x"4b"),
   414 => (x"ff",x"c3",x"48",x"d4"),
   415 => (x"bf",x"d0",x"ff",x"78"),
   416 => (x"c4",x"98",x"73",x"48"),
   417 => (x"98",x"70",x"58",x"a6"),
   418 => (x"ff",x"87",x"ce",x"02"),
   419 => (x"73",x"48",x"bf",x"d0"),
   420 => (x"58",x"a6",x"c4",x"98"),
   421 => (x"f2",x"05",x"98",x"70"),
   422 => (x"48",x"d0",x"ff",x"87"),
   423 => (x"ff",x"78",x"c3",x"c4"),
   424 => (x"ff",x"c3",x"48",x"d4"),
   425 => (x"c0",x"1e",x"72",x"78"),
   426 => (x"d1",x"c1",x"f0",x"ff"),
   427 => (x"87",x"f5",x"ed",x"49"),
   428 => (x"98",x"70",x"86",x"c4"),
   429 => (x"87",x"ee",x"c0",x"05"),
   430 => (x"d4",x"1e",x"c0",x"c8"),
   431 => (x"f8",x"fb",x"49",x"66"),
   432 => (x"70",x"86",x"c4",x"87"),
   433 => (x"bf",x"d0",x"ff",x"4c"),
   434 => (x"c4",x"98",x"73",x"48"),
   435 => (x"98",x"70",x"58",x"a6"),
   436 => (x"ff",x"87",x"ce",x"02"),
   437 => (x"73",x"48",x"bf",x"d0"),
   438 => (x"58",x"a6",x"c4",x"98"),
   439 => (x"f2",x"05",x"98",x"70"),
   440 => (x"48",x"d0",x"ff",x"87"),
   441 => (x"48",x"74",x"78",x"c2"),
   442 => (x"87",x"f3",x"ec",x"26"),
   443 => (x"5c",x"5b",x"5e",x"0e"),
   444 => (x"c0",x"1e",x"0e",x"5d"),
   445 => (x"f0",x"ff",x"c0",x"1e"),
   446 => (x"ec",x"49",x"c9",x"c1"),
   447 => (x"1e",x"d2",x"87",x"e7"),
   448 => (x"49",x"da",x"ec",x"c2"),
   449 => (x"c8",x"87",x"f2",x"fa"),
   450 => (x"c1",x"4d",x"c0",x"86"),
   451 => (x"ad",x"b7",x"d2",x"85"),
   452 => (x"c2",x"87",x"f8",x"04"),
   453 => (x"bf",x"97",x"da",x"ec"),
   454 => (x"99",x"c0",x"c3",x"49"),
   455 => (x"05",x"a9",x"c0",x"c1"),
   456 => (x"c2",x"87",x"e7",x"c0"),
   457 => (x"bf",x"97",x"e1",x"ec"),
   458 => (x"c2",x"31",x"d0",x"49"),
   459 => (x"bf",x"97",x"e2",x"ec"),
   460 => (x"72",x"32",x"c8",x"4a"),
   461 => (x"e3",x"ec",x"c2",x"b1"),
   462 => (x"b1",x"4a",x"bf",x"97"),
   463 => (x"ff",x"cf",x"4d",x"71"),
   464 => (x"c1",x"9d",x"ff",x"ff"),
   465 => (x"c2",x"35",x"ca",x"85"),
   466 => (x"ec",x"c2",x"87",x"de"),
   467 => (x"4b",x"bf",x"97",x"e3"),
   468 => (x"9b",x"c6",x"33",x"c1"),
   469 => (x"97",x"e4",x"ec",x"c2"),
   470 => (x"b7",x"c7",x"49",x"bf"),
   471 => (x"c2",x"b3",x"71",x"29"),
   472 => (x"bf",x"97",x"df",x"ec"),
   473 => (x"98",x"cf",x"48",x"49"),
   474 => (x"c2",x"58",x"a6",x"c4"),
   475 => (x"bf",x"97",x"e0",x"ec"),
   476 => (x"ca",x"9c",x"c3",x"4c"),
   477 => (x"e1",x"ec",x"c2",x"34"),
   478 => (x"c2",x"49",x"bf",x"97"),
   479 => (x"c2",x"b4",x"71",x"31"),
   480 => (x"bf",x"97",x"e2",x"ec"),
   481 => (x"99",x"c0",x"c3",x"49"),
   482 => (x"71",x"29",x"b7",x"c6"),
   483 => (x"70",x"1e",x"74",x"b4"),
   484 => (x"cf",x"1e",x"73",x"1e"),
   485 => (x"e3",x"e3",x"1e",x"c6"),
   486 => (x"c1",x"83",x"c2",x"87"),
   487 => (x"70",x"30",x"73",x"48"),
   488 => (x"f3",x"cf",x"1e",x"4b"),
   489 => (x"87",x"d4",x"e3",x"1e"),
   490 => (x"66",x"d8",x"48",x"c1"),
   491 => (x"58",x"a6",x"dc",x"30"),
   492 => (x"4d",x"49",x"a4",x"c1"),
   493 => (x"1e",x"70",x"95",x"73"),
   494 => (x"fc",x"cf",x"1e",x"75"),
   495 => (x"87",x"fc",x"e2",x"1e"),
   496 => (x"6e",x"86",x"e4",x"c0"),
   497 => (x"b7",x"c0",x"c8",x"48"),
   498 => (x"87",x"d2",x"06",x"a8"),
   499 => (x"48",x"6e",x"35",x"c1"),
   500 => (x"c4",x"28",x"b7",x"c1"),
   501 => (x"c0",x"c8",x"58",x"a6"),
   502 => (x"ff",x"01",x"a8",x"b7"),
   503 => (x"1e",x"75",x"87",x"ee"),
   504 => (x"e2",x"1e",x"d2",x"d0"),
   505 => (x"86",x"c8",x"87",x"d6"),
   506 => (x"e8",x"26",x"48",x"75"),
   507 => (x"5e",x"0e",x"87",x"ef"),
   508 => (x"71",x"0e",x"5c",x"5b"),
   509 => (x"d0",x"4c",x"c0",x"4b"),
   510 => (x"b7",x"c0",x"48",x"66"),
   511 => (x"e3",x"c0",x"06",x"a8"),
   512 => (x"cc",x"4a",x"13",x"87"),
   513 => (x"49",x"bf",x"97",x"66"),
   514 => (x"c1",x"48",x"66",x"cc"),
   515 => (x"58",x"a6",x"d0",x"80"),
   516 => (x"02",x"aa",x"b7",x"71"),
   517 => (x"48",x"c1",x"87",x"c4"),
   518 => (x"84",x"c1",x"87",x"cc"),
   519 => (x"ac",x"b7",x"66",x"d0"),
   520 => (x"87",x"dd",x"ff",x"04"),
   521 => (x"87",x"c2",x"48",x"c0"),
   522 => (x"4c",x"26",x"4d",x"26"),
   523 => (x"4f",x"26",x"4b",x"26"),
   524 => (x"5c",x"5b",x"5e",x"0e"),
   525 => (x"f5",x"c2",x"0e",x"5d"),
   526 => (x"78",x"c0",x"48",x"c0"),
   527 => (x"49",x"dd",x"ef",x"c0"),
   528 => (x"c2",x"87",x"e4",x"e5"),
   529 => (x"c0",x"1e",x"f8",x"ec"),
   530 => (x"87",x"dd",x"f8",x"49"),
   531 => (x"98",x"70",x"86",x"c4"),
   532 => (x"c0",x"87",x"cc",x"05"),
   533 => (x"e5",x"49",x"c9",x"ec"),
   534 => (x"48",x"c0",x"87",x"cd"),
   535 => (x"c0",x"87",x"e7",x"ca"),
   536 => (x"e5",x"49",x"ea",x"ef"),
   537 => (x"4b",x"c0",x"87",x"c1"),
   538 => (x"48",x"f8",x"f9",x"c2"),
   539 => (x"1e",x"c8",x"78",x"c1"),
   540 => (x"1e",x"c1",x"f0",x"c0"),
   541 => (x"49",x"ee",x"ed",x"c2"),
   542 => (x"c8",x"87",x"f3",x"fd"),
   543 => (x"05",x"98",x"70",x"86"),
   544 => (x"f9",x"c2",x"87",x"c6"),
   545 => (x"78",x"c0",x"48",x"f8"),
   546 => (x"f0",x"c0",x"1e",x"c8"),
   547 => (x"ee",x"c2",x"1e",x"ca"),
   548 => (x"d9",x"fd",x"49",x"ca"),
   549 => (x"70",x"86",x"c8",x"87"),
   550 => (x"87",x"c6",x"05",x"98"),
   551 => (x"48",x"f8",x"f9",x"c2"),
   552 => (x"f9",x"c2",x"78",x"c0"),
   553 => (x"c0",x"1e",x"bf",x"f8"),
   554 => (x"ff",x"1e",x"d3",x"f0"),
   555 => (x"c8",x"87",x"cd",x"df"),
   556 => (x"f8",x"f9",x"c2",x"86"),
   557 => (x"f7",x"c1",x"02",x"bf"),
   558 => (x"f6",x"f4",x"c2",x"87"),
   559 => (x"1e",x"49",x"bf",x"9f"),
   560 => (x"49",x"f6",x"f4",x"c2"),
   561 => (x"a0",x"c2",x"f8",x"48"),
   562 => (x"d0",x"1e",x"71",x"89"),
   563 => (x"1e",x"c0",x"c8",x"1e"),
   564 => (x"1e",x"fb",x"ec",x"c0"),
   565 => (x"87",x"e4",x"de",x"ff"),
   566 => (x"f3",x"c2",x"86",x"d4"),
   567 => (x"c2",x"4b",x"bf",x"fe"),
   568 => (x"bf",x"9f",x"f6",x"f4"),
   569 => (x"ea",x"d6",x"c5",x"4a"),
   570 => (x"c8",x"c0",x"05",x"aa"),
   571 => (x"fe",x"f3",x"c2",x"87"),
   572 => (x"d4",x"c0",x"4b",x"bf"),
   573 => (x"d5",x"e9",x"ca",x"87"),
   574 => (x"cc",x"c0",x"02",x"aa"),
   575 => (x"dd",x"ec",x"c0",x"87"),
   576 => (x"87",x"e3",x"e2",x"49"),
   577 => (x"fd",x"c7",x"48",x"c0"),
   578 => (x"c0",x"1e",x"73",x"87"),
   579 => (x"ff",x"1e",x"f8",x"ed"),
   580 => (x"c2",x"87",x"e9",x"dd"),
   581 => (x"73",x"1e",x"f8",x"ec"),
   582 => (x"87",x"cd",x"f5",x"49"),
   583 => (x"98",x"70",x"86",x"cc"),
   584 => (x"87",x"c5",x"c0",x"05"),
   585 => (x"dd",x"c7",x"48",x"c0"),
   586 => (x"d0",x"ee",x"c0",x"87"),
   587 => (x"87",x"f7",x"e1",x"49"),
   588 => (x"1e",x"e6",x"f0",x"c0"),
   589 => (x"87",x"c4",x"dd",x"ff"),
   590 => (x"f0",x"c0",x"1e",x"c8"),
   591 => (x"ee",x"c2",x"1e",x"fe"),
   592 => (x"e9",x"fa",x"49",x"ca"),
   593 => (x"70",x"86",x"cc",x"87"),
   594 => (x"c9",x"c0",x"05",x"98"),
   595 => (x"c0",x"f5",x"c2",x"87"),
   596 => (x"c0",x"78",x"c1",x"48"),
   597 => (x"1e",x"c8",x"87",x"e4"),
   598 => (x"1e",x"c7",x"f1",x"c0"),
   599 => (x"49",x"ee",x"ed",x"c2"),
   600 => (x"c8",x"87",x"cb",x"fa"),
   601 => (x"02",x"98",x"70",x"86"),
   602 => (x"c0",x"87",x"cf",x"c0"),
   603 => (x"ff",x"1e",x"f7",x"ee"),
   604 => (x"c4",x"87",x"c9",x"dc"),
   605 => (x"c6",x"48",x"c0",x"86"),
   606 => (x"f4",x"c2",x"87",x"cc"),
   607 => (x"49",x"bf",x"97",x"f6"),
   608 => (x"05",x"a9",x"d5",x"c1"),
   609 => (x"c2",x"87",x"cd",x"c0"),
   610 => (x"bf",x"97",x"f7",x"f4"),
   611 => (x"a9",x"ea",x"c2",x"49"),
   612 => (x"87",x"c5",x"c0",x"02"),
   613 => (x"ed",x"c5",x"48",x"c0"),
   614 => (x"f8",x"ec",x"c2",x"87"),
   615 => (x"c3",x"4c",x"bf",x"97"),
   616 => (x"c0",x"02",x"ac",x"e9"),
   617 => (x"eb",x"c3",x"87",x"cc"),
   618 => (x"c5",x"c0",x"02",x"ac"),
   619 => (x"c5",x"48",x"c0",x"87"),
   620 => (x"ed",x"c2",x"87",x"d4"),
   621 => (x"49",x"bf",x"97",x"c3"),
   622 => (x"cc",x"c0",x"05",x"99"),
   623 => (x"c4",x"ed",x"c2",x"87"),
   624 => (x"c2",x"49",x"bf",x"97"),
   625 => (x"c5",x"c0",x"02",x"a9"),
   626 => (x"c4",x"48",x"c0",x"87"),
   627 => (x"ed",x"c2",x"87",x"f8"),
   628 => (x"48",x"bf",x"97",x"c5"),
   629 => (x"58",x"fc",x"f4",x"c2"),
   630 => (x"c1",x"4a",x"49",x"70"),
   631 => (x"c0",x"f5",x"c2",x"8a"),
   632 => (x"71",x"1e",x"72",x"5a"),
   633 => (x"d0",x"f1",x"c0",x"1e"),
   634 => (x"cf",x"da",x"ff",x"1e"),
   635 => (x"c2",x"86",x"cc",x"87"),
   636 => (x"bf",x"97",x"c6",x"ed"),
   637 => (x"c2",x"81",x"73",x"49"),
   638 => (x"bf",x"97",x"c7",x"ed"),
   639 => (x"35",x"c8",x"4d",x"4a"),
   640 => (x"f9",x"c2",x"85",x"71"),
   641 => (x"ed",x"c2",x"5d",x"d8"),
   642 => (x"48",x"bf",x"97",x"c8"),
   643 => (x"58",x"ec",x"f9",x"c2"),
   644 => (x"bf",x"c0",x"f5",x"c2"),
   645 => (x"87",x"dc",x"c2",x"02"),
   646 => (x"ef",x"c0",x"1e",x"c8"),
   647 => (x"ee",x"c2",x"1e",x"d4"),
   648 => (x"c9",x"f7",x"49",x"ca"),
   649 => (x"70",x"86",x"c8",x"87"),
   650 => (x"c5",x"c0",x"02",x"98"),
   651 => (x"c3",x"48",x"c0",x"87"),
   652 => (x"f4",x"c2",x"87",x"d4"),
   653 => (x"48",x"4a",x"bf",x"f8"),
   654 => (x"f5",x"c2",x"30",x"c4"),
   655 => (x"f9",x"c2",x"58",x"c8"),
   656 => (x"ed",x"c2",x"5a",x"e8"),
   657 => (x"49",x"bf",x"97",x"dd"),
   658 => (x"ed",x"c2",x"31",x"c8"),
   659 => (x"4b",x"bf",x"97",x"dc"),
   660 => (x"ed",x"c2",x"49",x"a1"),
   661 => (x"4b",x"bf",x"97",x"de"),
   662 => (x"a1",x"73",x"33",x"d0"),
   663 => (x"df",x"ed",x"c2",x"49"),
   664 => (x"d8",x"4b",x"bf",x"97"),
   665 => (x"49",x"a1",x"73",x"33"),
   666 => (x"59",x"f0",x"f9",x"c2"),
   667 => (x"bf",x"e8",x"f9",x"c2"),
   668 => (x"d4",x"f9",x"c2",x"91"),
   669 => (x"f9",x"c2",x"81",x"bf"),
   670 => (x"ed",x"c2",x"59",x"dc"),
   671 => (x"4b",x"bf",x"97",x"e5"),
   672 => (x"ed",x"c2",x"33",x"c8"),
   673 => (x"4c",x"bf",x"97",x"e4"),
   674 => (x"ed",x"c2",x"4b",x"a3"),
   675 => (x"4c",x"bf",x"97",x"e6"),
   676 => (x"a3",x"74",x"34",x"d0"),
   677 => (x"e7",x"ed",x"c2",x"4b"),
   678 => (x"cf",x"4c",x"bf",x"97"),
   679 => (x"74",x"34",x"d8",x"9c"),
   680 => (x"f9",x"c2",x"4b",x"a3"),
   681 => (x"8b",x"c2",x"5b",x"e0"),
   682 => (x"f9",x"c2",x"92",x"73"),
   683 => (x"a1",x"72",x"48",x"e0"),
   684 => (x"87",x"cb",x"c1",x"78"),
   685 => (x"97",x"ca",x"ed",x"c2"),
   686 => (x"31",x"c8",x"49",x"bf"),
   687 => (x"97",x"c9",x"ed",x"c2"),
   688 => (x"49",x"a1",x"4a",x"bf"),
   689 => (x"59",x"c8",x"f5",x"c2"),
   690 => (x"ff",x"c7",x"31",x"c5"),
   691 => (x"c2",x"29",x"c9",x"81"),
   692 => (x"c2",x"59",x"e8",x"f9"),
   693 => (x"bf",x"97",x"cf",x"ed"),
   694 => (x"c2",x"32",x"c8",x"4a"),
   695 => (x"bf",x"97",x"ce",x"ed"),
   696 => (x"c2",x"4a",x"a2",x"4b"),
   697 => (x"c2",x"5a",x"f0",x"f9"),
   698 => (x"92",x"bf",x"e8",x"f9"),
   699 => (x"f9",x"c2",x"82",x"75"),
   700 => (x"f9",x"c2",x"5a",x"e4"),
   701 => (x"78",x"c0",x"48",x"dc"),
   702 => (x"48",x"d8",x"f9",x"c2"),
   703 => (x"c0",x"78",x"a1",x"72"),
   704 => (x"87",x"e3",x"cd",x"49"),
   705 => (x"df",x"f4",x"48",x"c1"),
   706 => (x"61",x"65",x"52",x"87"),
   707 => (x"66",x"6f",x"20",x"64"),
   708 => (x"52",x"42",x"4d",x"20"),
   709 => (x"69",x"61",x"66",x"20"),
   710 => (x"0a",x"64",x"65",x"6c"),
   711 => (x"20",x"6f",x"4e",x"00"),
   712 => (x"74",x"72",x"61",x"70"),
   713 => (x"6f",x"69",x"74",x"69"),
   714 => (x"69",x"73",x"20",x"6e"),
   715 => (x"74",x"61",x"6e",x"67"),
   716 => (x"20",x"65",x"72",x"75"),
   717 => (x"6e",x"75",x"6f",x"66"),
   718 => (x"4d",x"00",x"0a",x"64"),
   719 => (x"69",x"73",x"52",x"42"),
   720 => (x"20",x"3a",x"65",x"7a"),
   721 => (x"20",x"2c",x"64",x"25"),
   722 => (x"74",x"72",x"61",x"70"),
   723 => (x"6f",x"69",x"74",x"69"),
   724 => (x"7a",x"69",x"73",x"6e"),
   725 => (x"25",x"20",x"3a",x"65"),
   726 => (x"6f",x"20",x"2c",x"64"),
   727 => (x"65",x"73",x"66",x"66"),
   728 => (x"66",x"6f",x"20",x"74"),
   729 => (x"67",x"69",x"73",x"20"),
   730 => (x"64",x"25",x"20",x"3a"),
   731 => (x"69",x"73",x"20",x"2c"),
   732 => (x"78",x"30",x"20",x"67"),
   733 => (x"00",x"0a",x"78",x"25"),
   734 => (x"64",x"61",x"65",x"52"),
   735 => (x"20",x"67",x"6e",x"69"),
   736 => (x"74",x"6f",x"6f",x"62"),
   737 => (x"63",x"65",x"73",x"20"),
   738 => (x"20",x"72",x"6f",x"74"),
   739 => (x"00",x"0a",x"64",x"25"),
   740 => (x"64",x"61",x"65",x"52"),
   741 => (x"6f",x"6f",x"62",x"20"),
   742 => (x"65",x"73",x"20",x"74"),
   743 => (x"72",x"6f",x"74",x"63"),
   744 => (x"6f",x"72",x"66",x"20"),
   745 => (x"69",x"66",x"20",x"6d"),
   746 => (x"20",x"74",x"73",x"72"),
   747 => (x"74",x"72",x"61",x"70"),
   748 => (x"6f",x"69",x"74",x"69"),
   749 => (x"55",x"00",x"0a",x"6e"),
   750 => (x"70",x"75",x"73",x"6e"),
   751 => (x"74",x"72",x"6f",x"70"),
   752 => (x"70",x"20",x"64",x"65"),
   753 => (x"69",x"74",x"72",x"61"),
   754 => (x"6e",x"6f",x"69",x"74"),
   755 => (x"70",x"79",x"74",x"20"),
   756 => (x"00",x"0d",x"21",x"65"),
   757 => (x"33",x"54",x"41",x"46"),
   758 => (x"20",x"20",x"20",x"32"),
   759 => (x"61",x"65",x"52",x"00"),
   760 => (x"67",x"6e",x"69",x"64"),
   761 => (x"52",x"42",x"4d",x"20"),
   762 => (x"42",x"4d",x"00",x"0a"),
   763 => (x"75",x"73",x"20",x"52"),
   764 => (x"73",x"65",x"63",x"63"),
   765 => (x"6c",x"75",x"66",x"73"),
   766 => (x"72",x"20",x"79",x"6c"),
   767 => (x"0a",x"64",x"61",x"65"),
   768 => (x"54",x"41",x"46",x"00"),
   769 => (x"20",x"20",x"36",x"31"),
   770 => (x"41",x"46",x"00",x"20"),
   771 => (x"20",x"32",x"33",x"54"),
   772 => (x"50",x"00",x"20",x"20"),
   773 => (x"69",x"74",x"72",x"61"),
   774 => (x"6e",x"6f",x"69",x"74"),
   775 => (x"6e",x"75",x"6f",x"63"),
   776 => (x"64",x"25",x"20",x"74"),
   777 => (x"75",x"48",x"00",x"0a"),
   778 => (x"6e",x"69",x"74",x"6e"),
   779 => (x"6f",x"66",x"20",x"67"),
   780 => (x"69",x"66",x"20",x"72"),
   781 => (x"79",x"73",x"65",x"6c"),
   782 => (x"6d",x"65",x"74",x"73"),
   783 => (x"41",x"46",x"00",x"0a"),
   784 => (x"20",x"32",x"33",x"54"),
   785 => (x"46",x"00",x"20",x"20"),
   786 => (x"36",x"31",x"54",x"41"),
   787 => (x"00",x"20",x"20",x"20"),
   788 => (x"73",x"75",x"6c",x"43"),
   789 => (x"20",x"72",x"65",x"74"),
   790 => (x"65",x"7a",x"69",x"73"),
   791 => (x"64",x"25",x"20",x"3a"),
   792 => (x"6c",x"43",x"20",x"2c"),
   793 => (x"65",x"74",x"73",x"75"),
   794 => (x"61",x"6d",x"20",x"72"),
   795 => (x"20",x"2c",x"6b",x"73"),
   796 => (x"00",x"0a",x"64",x"25"),
   797 => (x"6e",x"65",x"70",x"4f"),
   798 => (x"66",x"20",x"64",x"65"),
   799 => (x"2c",x"65",x"6c",x"69"),
   800 => (x"61",x"6f",x"6c",x"20"),
   801 => (x"67",x"6e",x"69",x"64"),
   802 => (x"0a",x"2e",x"2e",x"2e"),
   803 => (x"6e",x"61",x"43",x"00"),
   804 => (x"6f",x"20",x"74",x"27"),
   805 => (x"20",x"6e",x"65",x"70"),
   806 => (x"00",x"0a",x"73",x"25"),
   807 => (x"5c",x"5b",x"5e",x"0e"),
   808 => (x"4a",x"71",x"0e",x"5d"),
   809 => (x"bf",x"c0",x"f5",x"c2"),
   810 => (x"72",x"87",x"cc",x"02"),
   811 => (x"2b",x"b7",x"c7",x"4b"),
   812 => (x"ff",x"c1",x"4d",x"72"),
   813 => (x"72",x"87",x"ca",x"9d"),
   814 => (x"2b",x"b7",x"c8",x"4b"),
   815 => (x"ff",x"c3",x"4d",x"72"),
   816 => (x"f8",x"ec",x"c2",x"9d"),
   817 => (x"d4",x"f9",x"c2",x"1e"),
   818 => (x"81",x"73",x"49",x"bf"),
   819 => (x"87",x"d9",x"e6",x"71"),
   820 => (x"98",x"70",x"86",x"c4"),
   821 => (x"c0",x"87",x"c5",x"05"),
   822 => (x"87",x"e6",x"c0",x"48"),
   823 => (x"bf",x"c0",x"f5",x"c2"),
   824 => (x"75",x"87",x"d2",x"02"),
   825 => (x"c2",x"91",x"c4",x"49"),
   826 => (x"69",x"81",x"f8",x"ec"),
   827 => (x"ff",x"ff",x"cf",x"4c"),
   828 => (x"cb",x"9c",x"ff",x"ff"),
   829 => (x"c2",x"49",x"75",x"87"),
   830 => (x"f8",x"ec",x"c2",x"91"),
   831 => (x"4c",x"69",x"9f",x"81"),
   832 => (x"e3",x"ec",x"48",x"74"),
   833 => (x"5b",x"5e",x"0e",x"87"),
   834 => (x"f4",x"0e",x"5d",x"5c"),
   835 => (x"c0",x"4c",x"71",x"86"),
   836 => (x"f0",x"f9",x"c2",x"4b"),
   837 => (x"a6",x"c4",x"7e",x"bf"),
   838 => (x"f4",x"f9",x"c2",x"48"),
   839 => (x"a6",x"c8",x"78",x"bf"),
   840 => (x"c2",x"78",x"c0",x"48"),
   841 => (x"48",x"bf",x"c4",x"f5"),
   842 => (x"c2",x"06",x"a8",x"c0"),
   843 => (x"66",x"c8",x"87",x"e3"),
   844 => (x"05",x"99",x"cf",x"49"),
   845 => (x"ec",x"c2",x"87",x"d8"),
   846 => (x"66",x"c8",x"1e",x"f8"),
   847 => (x"80",x"c1",x"48",x"49"),
   848 => (x"e4",x"58",x"a6",x"cc"),
   849 => (x"86",x"c4",x"87",x"e3"),
   850 => (x"4b",x"f8",x"ec",x"c2"),
   851 => (x"e0",x"c0",x"87",x"c3"),
   852 => (x"4a",x"6b",x"97",x"83"),
   853 => (x"e7",x"c1",x"02",x"9a"),
   854 => (x"aa",x"e5",x"c3",x"87"),
   855 => (x"87",x"e0",x"c1",x"02"),
   856 => (x"97",x"49",x"a3",x"cb"),
   857 => (x"99",x"d8",x"49",x"69"),
   858 => (x"87",x"d4",x"c1",x"05"),
   859 => (x"d0",x"ff",x"49",x"73"),
   860 => (x"1e",x"cb",x"87",x"f5"),
   861 => (x"1e",x"66",x"e0",x"c0"),
   862 => (x"f1",x"e9",x"49",x"73"),
   863 => (x"70",x"86",x"c8",x"87"),
   864 => (x"fb",x"c0",x"05",x"98"),
   865 => (x"4a",x"a3",x"dc",x"87"),
   866 => (x"6a",x"49",x"a4",x"c4"),
   867 => (x"49",x"a3",x"da",x"79"),
   868 => (x"9f",x"4d",x"a4",x"c8"),
   869 => (x"c2",x"7d",x"48",x"69"),
   870 => (x"02",x"bf",x"c0",x"f5"),
   871 => (x"a3",x"d4",x"87",x"d3"),
   872 => (x"49",x"69",x"9f",x"49"),
   873 => (x"99",x"ff",x"ff",x"c0"),
   874 => (x"30",x"d0",x"48",x"71"),
   875 => (x"c2",x"58",x"a6",x"c4"),
   876 => (x"6e",x"7e",x"c0",x"87"),
   877 => (x"70",x"80",x"6d",x"48"),
   878 => (x"c1",x"7c",x"c0",x"7d"),
   879 => (x"87",x"c5",x"c1",x"48"),
   880 => (x"c1",x"48",x"66",x"c8"),
   881 => (x"58",x"a6",x"cc",x"80"),
   882 => (x"bf",x"c4",x"f5",x"c2"),
   883 => (x"dd",x"fd",x"04",x"a8"),
   884 => (x"c0",x"f5",x"c2",x"87"),
   885 => (x"ea",x"c0",x"02",x"bf"),
   886 => (x"fa",x"49",x"6e",x"87"),
   887 => (x"a6",x"c4",x"87",x"fe"),
   888 => (x"cf",x"49",x"70",x"58"),
   889 => (x"f8",x"ff",x"ff",x"ff"),
   890 => (x"d6",x"02",x"a9",x"99"),
   891 => (x"c2",x"49",x"70",x"87"),
   892 => (x"f8",x"f4",x"c2",x"89"),
   893 => (x"f9",x"c2",x"91",x"bf"),
   894 => (x"71",x"48",x"bf",x"d8"),
   895 => (x"58",x"a6",x"c8",x"80"),
   896 => (x"c0",x"87",x"db",x"fc"),
   897 => (x"e8",x"8e",x"f4",x"48"),
   898 => (x"73",x"1e",x"87",x"de"),
   899 => (x"6a",x"4a",x"71",x"1e"),
   900 => (x"71",x"81",x"c1",x"49"),
   901 => (x"fc",x"f4",x"c2",x"7a"),
   902 => (x"cb",x"05",x"99",x"bf"),
   903 => (x"4b",x"a2",x"c8",x"87"),
   904 => (x"f7",x"f9",x"49",x"6b"),
   905 => (x"7b",x"49",x"70",x"87"),
   906 => (x"ff",x"e7",x"48",x"c1"),
   907 => (x"1e",x"73",x"1e",x"87"),
   908 => (x"f9",x"c2",x"4b",x"71"),
   909 => (x"c8",x"49",x"bf",x"d8"),
   910 => (x"4a",x"6a",x"4a",x"a3"),
   911 => (x"f4",x"c2",x"8a",x"c2"),
   912 => (x"72",x"92",x"bf",x"f8"),
   913 => (x"f4",x"c2",x"49",x"a1"),
   914 => (x"6b",x"4a",x"bf",x"fc"),
   915 => (x"49",x"a1",x"72",x"9a"),
   916 => (x"71",x"1e",x"66",x"c8"),
   917 => (x"c4",x"87",x"d2",x"e0"),
   918 => (x"05",x"98",x"70",x"86"),
   919 => (x"48",x"c0",x"87",x"c4"),
   920 => (x"48",x"c1",x"87",x"c2"),
   921 => (x"0e",x"87",x"c5",x"e7"),
   922 => (x"0e",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"c0",x"4a",x"71"),
   924 => (x"c0",x"02",x"9a",x"72"),
   925 => (x"a2",x"da",x"87",x"e0"),
   926 => (x"4b",x"69",x"9f",x"49"),
   927 => (x"bf",x"c0",x"f5",x"c2"),
   928 => (x"d4",x"87",x"cf",x"02"),
   929 => (x"69",x"9f",x"49",x"a2"),
   930 => (x"ff",x"c0",x"4c",x"49"),
   931 => (x"34",x"d0",x"9c",x"ff"),
   932 => (x"4c",x"c0",x"87",x"c2"),
   933 => (x"9b",x"73",x"b3",x"74"),
   934 => (x"4a",x"87",x"df",x"02"),
   935 => (x"f4",x"c2",x"8a",x"c2"),
   936 => (x"92",x"49",x"bf",x"f8"),
   937 => (x"bf",x"d8",x"f9",x"c2"),
   938 => (x"c2",x"80",x"72",x"48"),
   939 => (x"71",x"58",x"f8",x"f9"),
   940 => (x"c2",x"30",x"c4",x"48"),
   941 => (x"c0",x"58",x"c8",x"f5"),
   942 => (x"f9",x"c2",x"87",x"e9"),
   943 => (x"c2",x"4b",x"bf",x"dc"),
   944 => (x"c2",x"48",x"f4",x"f9"),
   945 => (x"78",x"bf",x"e0",x"f9"),
   946 => (x"bf",x"c0",x"f5",x"c2"),
   947 => (x"c2",x"87",x"c9",x"02"),
   948 => (x"49",x"bf",x"f8",x"f4"),
   949 => (x"87",x"c7",x"31",x"c4"),
   950 => (x"bf",x"e4",x"f9",x"c2"),
   951 => (x"c2",x"31",x"c4",x"49"),
   952 => (x"c2",x"59",x"c8",x"f5"),
   953 => (x"e5",x"5b",x"f4",x"f9"),
   954 => (x"5e",x"0e",x"87",x"c0"),
   955 => (x"0e",x"5d",x"5c",x"5b"),
   956 => (x"9a",x"4a",x"71",x"1e"),
   957 => (x"c2",x"87",x"de",x"02"),
   958 => (x"c0",x"48",x"f4",x"ec"),
   959 => (x"ec",x"ec",x"c2",x"78"),
   960 => (x"f4",x"f9",x"c2",x"48"),
   961 => (x"ec",x"c2",x"78",x"bf"),
   962 => (x"f9",x"c2",x"48",x"f0"),
   963 => (x"c1",x"78",x"bf",x"f0"),
   964 => (x"c0",x"48",x"e2",x"c2"),
   965 => (x"c4",x"f5",x"c2",x"78"),
   966 => (x"ec",x"c2",x"49",x"bf"),
   967 => (x"71",x"4a",x"bf",x"f4"),
   968 => (x"fe",x"c3",x"03",x"aa"),
   969 => (x"cf",x"49",x"72",x"87"),
   970 => (x"e1",x"c0",x"05",x"99"),
   971 => (x"f8",x"ec",x"c2",x"87"),
   972 => (x"ec",x"ec",x"c2",x"1e"),
   973 => (x"ec",x"c2",x"49",x"bf"),
   974 => (x"a1",x"c1",x"48",x"ec"),
   975 => (x"dc",x"ff",x"71",x"78"),
   976 => (x"86",x"c4",x"87",x"e7"),
   977 => (x"48",x"de",x"c2",x"c1"),
   978 => (x"78",x"f8",x"ec",x"c2"),
   979 => (x"c2",x"c1",x"87",x"cc"),
   980 => (x"c0",x"48",x"bf",x"de"),
   981 => (x"c2",x"c1",x"80",x"e0"),
   982 => (x"ec",x"c2",x"58",x"e2"),
   983 => (x"c1",x"48",x"bf",x"f4"),
   984 => (x"f8",x"ec",x"c2",x"80"),
   985 => (x"de",x"c2",x"c1",x"58"),
   986 => (x"a3",x"cb",x"4b",x"bf"),
   987 => (x"cf",x"4c",x"11",x"49"),
   988 => (x"dd",x"c1",x"05",x"ac"),
   989 => (x"10",x"9e",x"27",x"87"),
   990 => (x"97",x"bf",x"00",x"00"),
   991 => (x"99",x"df",x"49",x"bf"),
   992 => (x"91",x"cd",x"89",x"c1"),
   993 => (x"81",x"c8",x"f5",x"c2"),
   994 => (x"12",x"4a",x"a3",x"c1"),
   995 => (x"4a",x"a3",x"c3",x"51"),
   996 => (x"a3",x"c5",x"51",x"12"),
   997 => (x"c7",x"51",x"12",x"4a"),
   998 => (x"51",x"12",x"4a",x"a3"),
   999 => (x"12",x"4a",x"a3",x"c9"),
  1000 => (x"4a",x"a3",x"ce",x"51"),
  1001 => (x"a3",x"d0",x"51",x"12"),
  1002 => (x"d2",x"51",x"12",x"4a"),
  1003 => (x"51",x"12",x"4a",x"a3"),
  1004 => (x"12",x"4a",x"a3",x"d4"),
  1005 => (x"4a",x"a3",x"d6",x"51"),
  1006 => (x"a3",x"d8",x"51",x"12"),
  1007 => (x"dc",x"51",x"12",x"4a"),
  1008 => (x"51",x"12",x"4a",x"a3"),
  1009 => (x"12",x"4a",x"a3",x"de"),
  1010 => (x"e2",x"c2",x"c1",x"51"),
  1011 => (x"c1",x"78",x"c1",x"48"),
  1012 => (x"49",x"74",x"87",x"c1"),
  1013 => (x"c0",x"05",x"99",x"c8"),
  1014 => (x"49",x"74",x"87",x"f3"),
  1015 => (x"d0",x"05",x"99",x"d0"),
  1016 => (x"02",x"66",x"d4",x"87"),
  1017 => (x"73",x"87",x"ca",x"c0"),
  1018 => (x"0f",x"66",x"d4",x"49"),
  1019 => (x"dc",x"02",x"98",x"70"),
  1020 => (x"e2",x"c2",x"c1",x"87"),
  1021 => (x"c6",x"c0",x"05",x"bf"),
  1022 => (x"c8",x"f5",x"c2",x"87"),
  1023 => (x"c1",x"50",x"c0",x"48"),
  1024 => (x"c0",x"48",x"e2",x"c2"),
  1025 => (x"de",x"c2",x"c1",x"78"),
  1026 => (x"cc",x"c2",x"48",x"bf"),
  1027 => (x"e2",x"c2",x"c1",x"87"),
  1028 => (x"c2",x"78",x"c0",x"48"),
  1029 => (x"49",x"bf",x"c4",x"f5"),
  1030 => (x"bf",x"f4",x"ec",x"c2"),
  1031 => (x"04",x"aa",x"71",x"4a"),
  1032 => (x"c2",x"87",x"c2",x"fc"),
  1033 => (x"05",x"bf",x"f4",x"f9"),
  1034 => (x"c2",x"87",x"c8",x"c0"),
  1035 => (x"02",x"bf",x"c0",x"f5"),
  1036 => (x"c2",x"87",x"e4",x"c1"),
  1037 => (x"49",x"bf",x"f0",x"ec"),
  1038 => (x"c2",x"87",x"e1",x"f1"),
  1039 => (x"70",x"58",x"f4",x"ec"),
  1040 => (x"c0",x"f5",x"c2",x"4d"),
  1041 => (x"d7",x"c0",x"02",x"bf"),
  1042 => (x"cf",x"49",x"75",x"87"),
  1043 => (x"f8",x"ff",x"ff",x"ff"),
  1044 => (x"c0",x"02",x"a9",x"99"),
  1045 => (x"4c",x"c0",x"87",x"c5"),
  1046 => (x"c1",x"87",x"d9",x"c0"),
  1047 => (x"87",x"d4",x"c0",x"4c"),
  1048 => (x"ff",x"cf",x"49",x"75"),
  1049 => (x"02",x"a9",x"99",x"f8"),
  1050 => (x"c0",x"87",x"c5",x"c0"),
  1051 => (x"87",x"c2",x"c0",x"7e"),
  1052 => (x"4c",x"6e",x"7e",x"c1"),
  1053 => (x"c0",x"05",x"9c",x"74"),
  1054 => (x"49",x"75",x"87",x"dd"),
  1055 => (x"f4",x"c2",x"89",x"c2"),
  1056 => (x"c2",x"91",x"bf",x"f8"),
  1057 => (x"48",x"bf",x"d8",x"f9"),
  1058 => (x"ec",x"c2",x"80",x"71"),
  1059 => (x"ec",x"c2",x"58",x"f0"),
  1060 => (x"78",x"c0",x"48",x"f4"),
  1061 => (x"c0",x"87",x"fe",x"f9"),
  1062 => (x"de",x"ff",x"26",x"48"),
  1063 => (x"00",x"00",x"87",x"ca"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"ff",x"1e",x"00",x"00"),
  1066 => (x"ff",x"c3",x"48",x"d4"),
  1067 => (x"99",x"49",x"68",x"78"),
  1068 => (x"c0",x"87",x"c6",x"02"),
  1069 => (x"ee",x"05",x"a9",x"fb"),
  1070 => (x"26",x"48",x"71",x"87"),
  1071 => (x"5b",x"5e",x"0e",x"4f"),
  1072 => (x"4a",x"71",x"0e",x"5c"),
  1073 => (x"d4",x"ff",x"4b",x"c0"),
  1074 => (x"78",x"ff",x"c3",x"48"),
  1075 => (x"02",x"99",x"49",x"68"),
  1076 => (x"c0",x"87",x"c1",x"c1"),
  1077 => (x"c0",x"02",x"a9",x"ec"),
  1078 => (x"fb",x"c0",x"87",x"fa"),
  1079 => (x"f3",x"c0",x"02",x"a9"),
  1080 => (x"b7",x"66",x"cc",x"87"),
  1081 => (x"87",x"cc",x"03",x"ab"),
  1082 => (x"c7",x"02",x"66",x"d0"),
  1083 => (x"97",x"09",x"72",x"87"),
  1084 => (x"82",x"c1",x"09",x"79"),
  1085 => (x"c2",x"02",x"99",x"71"),
  1086 => (x"ff",x"83",x"c1",x"87"),
  1087 => (x"ff",x"c3",x"48",x"d4"),
  1088 => (x"99",x"49",x"68",x"78"),
  1089 => (x"c0",x"87",x"cd",x"02"),
  1090 => (x"c7",x"02",x"a9",x"ec"),
  1091 => (x"a9",x"fb",x"c0",x"87"),
  1092 => (x"87",x"cd",x"ff",x"05"),
  1093 => (x"c3",x"02",x"66",x"d0"),
  1094 => (x"7a",x"97",x"c0",x"87"),
  1095 => (x"05",x"a9",x"fb",x"c0"),
  1096 => (x"4c",x"73",x"87",x"c7"),
  1097 => (x"c2",x"8c",x"0c",x"c0"),
  1098 => (x"74",x"4c",x"73",x"87"),
  1099 => (x"26",x"87",x"c2",x"48"),
  1100 => (x"26",x"4c",x"26",x"4d"),
  1101 => (x"1e",x"4f",x"26",x"4b"),
  1102 => (x"c3",x"48",x"d4",x"ff"),
  1103 => (x"49",x"68",x"78",x"ff"),
  1104 => (x"a9",x"b7",x"f0",x"c0"),
  1105 => (x"c0",x"87",x"ca",x"04"),
  1106 => (x"01",x"a9",x"b7",x"f9"),
  1107 => (x"f0",x"c0",x"87",x"c3"),
  1108 => (x"b7",x"c1",x"c1",x"89"),
  1109 => (x"87",x"ca",x"04",x"a9"),
  1110 => (x"a9",x"b7",x"c6",x"c1"),
  1111 => (x"c0",x"87",x"c3",x"01"),
  1112 => (x"48",x"71",x"89",x"f7"),
  1113 => (x"5e",x"0e",x"4f",x"26"),
  1114 => (x"0e",x"5d",x"5c",x"5b"),
  1115 => (x"4c",x"71",x"86",x"f4"),
  1116 => (x"c0",x"4b",x"d4",x"ff"),
  1117 => (x"ff",x"c3",x"7e",x"4d"),
  1118 => (x"bf",x"d0",x"ff",x"7b"),
  1119 => (x"c0",x"c0",x"c8",x"48"),
  1120 => (x"58",x"a6",x"c8",x"98"),
  1121 => (x"d0",x"02",x"98",x"70"),
  1122 => (x"bf",x"d0",x"ff",x"87"),
  1123 => (x"c0",x"c0",x"c8",x"48"),
  1124 => (x"58",x"a6",x"c8",x"98"),
  1125 => (x"f0",x"05",x"98",x"70"),
  1126 => (x"48",x"d0",x"ff",x"87"),
  1127 => (x"d4",x"78",x"e1",x"c0"),
  1128 => (x"87",x"c2",x"fc",x"7b"),
  1129 => (x"02",x"99",x"49",x"70"),
  1130 => (x"c3",x"87",x"c7",x"c1"),
  1131 => (x"a6",x"c8",x"7b",x"ff"),
  1132 => (x"c8",x"78",x"6b",x"48"),
  1133 => (x"fb",x"c0",x"48",x"66"),
  1134 => (x"87",x"c8",x"02",x"a8"),
  1135 => (x"bf",x"d0",x"fa",x"c2"),
  1136 => (x"87",x"ee",x"c0",x"02"),
  1137 => (x"99",x"71",x"4d",x"c1"),
  1138 => (x"87",x"e6",x"c0",x"02"),
  1139 => (x"02",x"a9",x"fb",x"c0"),
  1140 => (x"d1",x"fb",x"87",x"c3"),
  1141 => (x"7b",x"ff",x"c3",x"87"),
  1142 => (x"c6",x"c1",x"49",x"6b"),
  1143 => (x"87",x"cc",x"05",x"a9"),
  1144 => (x"7b",x"7b",x"ff",x"c3"),
  1145 => (x"6b",x"48",x"a6",x"c8"),
  1146 => (x"4d",x"49",x"c0",x"78"),
  1147 => (x"ff",x"05",x"99",x"71"),
  1148 => (x"9d",x"75",x"87",x"da"),
  1149 => (x"87",x"de",x"c1",x"05"),
  1150 => (x"6b",x"7b",x"ff",x"c3"),
  1151 => (x"7b",x"ff",x"c3",x"4a"),
  1152 => (x"6b",x"48",x"a6",x"c4"),
  1153 => (x"c1",x"48",x"6e",x"78"),
  1154 => (x"58",x"a6",x"c4",x"80"),
  1155 => (x"97",x"49",x"a4",x"c8"),
  1156 => (x"66",x"c8",x"49",x"69"),
  1157 => (x"87",x"da",x"05",x"a9"),
  1158 => (x"97",x"49",x"a4",x"c9"),
  1159 => (x"05",x"aa",x"49",x"69"),
  1160 => (x"a4",x"ca",x"87",x"d0"),
  1161 => (x"49",x"69",x"97",x"49"),
  1162 => (x"05",x"a9",x"66",x"c4"),
  1163 => (x"4d",x"c1",x"87",x"c4"),
  1164 => (x"66",x"c8",x"87",x"d6"),
  1165 => (x"a8",x"ec",x"c0",x"48"),
  1166 => (x"c8",x"87",x"c9",x"02"),
  1167 => (x"fb",x"c0",x"48",x"66"),
  1168 => (x"87",x"c4",x"05",x"a8"),
  1169 => (x"4d",x"c1",x"7e",x"c0"),
  1170 => (x"c8",x"7b",x"ff",x"c3"),
  1171 => (x"78",x"6b",x"48",x"a6"),
  1172 => (x"fe",x"02",x"9d",x"75"),
  1173 => (x"d0",x"ff",x"87",x"e2"),
  1174 => (x"c0",x"c8",x"48",x"bf"),
  1175 => (x"a6",x"c8",x"98",x"c0"),
  1176 => (x"02",x"98",x"70",x"58"),
  1177 => (x"d0",x"ff",x"87",x"d0"),
  1178 => (x"c0",x"c8",x"48",x"bf"),
  1179 => (x"a6",x"c8",x"98",x"c0"),
  1180 => (x"05",x"98",x"70",x"58"),
  1181 => (x"d0",x"ff",x"87",x"f0"),
  1182 => (x"78",x"e0",x"c0",x"48"),
  1183 => (x"8e",x"f4",x"48",x"6e"),
  1184 => (x"0e",x"87",x"ec",x"fa"),
  1185 => (x"5d",x"5c",x"5b",x"5e"),
  1186 => (x"c4",x"86",x"f4",x"0e"),
  1187 => (x"d0",x"ff",x"59",x"a6"),
  1188 => (x"c0",x"c0",x"c8",x"4c"),
  1189 => (x"c2",x"1e",x"6e",x"4b"),
  1190 => (x"e9",x"49",x"d4",x"fa"),
  1191 => (x"86",x"c4",x"87",x"e7"),
  1192 => (x"c6",x"02",x"98",x"70"),
  1193 => (x"fa",x"c2",x"87",x"cb"),
  1194 => (x"6e",x"4d",x"bf",x"d8"),
  1195 => (x"87",x"f6",x"fa",x"49"),
  1196 => (x"70",x"58",x"a6",x"c8"),
  1197 => (x"49",x"66",x"c4",x"1e"),
  1198 => (x"1e",x"71",x"81",x"c8"),
  1199 => (x"1e",x"f8",x"d0",x"c1"),
  1200 => (x"87",x"f8",x"f6",x"fe"),
  1201 => (x"48",x"6c",x"86",x"cc"),
  1202 => (x"a6",x"cc",x"98",x"73"),
  1203 => (x"02",x"98",x"70",x"58"),
  1204 => (x"48",x"6c",x"87",x"cc"),
  1205 => (x"a6",x"c4",x"98",x"73"),
  1206 => (x"05",x"98",x"70",x"58"),
  1207 => (x"7c",x"c5",x"87",x"f4"),
  1208 => (x"c1",x"48",x"d4",x"ff"),
  1209 => (x"fa",x"c2",x"78",x"d5"),
  1210 => (x"c1",x"49",x"bf",x"d0"),
  1211 => (x"4a",x"66",x"c4",x"81"),
  1212 => (x"32",x"c6",x"8a",x"c1"),
  1213 => (x"b0",x"71",x"48",x"72"),
  1214 => (x"78",x"08",x"d4",x"ff"),
  1215 => (x"98",x"73",x"48",x"6c"),
  1216 => (x"70",x"58",x"a6",x"c4"),
  1217 => (x"87",x"cc",x"02",x"98"),
  1218 => (x"98",x"73",x"48",x"6c"),
  1219 => (x"70",x"58",x"a6",x"c4"),
  1220 => (x"87",x"f4",x"05",x"98"),
  1221 => (x"d4",x"ff",x"7c",x"c4"),
  1222 => (x"78",x"ff",x"c3",x"48"),
  1223 => (x"98",x"73",x"48",x"6c"),
  1224 => (x"70",x"58",x"a6",x"c4"),
  1225 => (x"87",x"cc",x"02",x"98"),
  1226 => (x"98",x"73",x"48",x"6c"),
  1227 => (x"70",x"58",x"a6",x"c4"),
  1228 => (x"87",x"f4",x"05",x"98"),
  1229 => (x"d4",x"ff",x"7c",x"c5"),
  1230 => (x"78",x"d3",x"c1",x"48"),
  1231 => (x"48",x"6c",x"78",x"c1"),
  1232 => (x"a6",x"c4",x"98",x"73"),
  1233 => (x"02",x"98",x"70",x"58"),
  1234 => (x"48",x"6c",x"87",x"cc"),
  1235 => (x"a6",x"c4",x"98",x"73"),
  1236 => (x"05",x"98",x"70",x"58"),
  1237 => (x"7c",x"c4",x"87",x"f4"),
  1238 => (x"c2",x"02",x"9d",x"75"),
  1239 => (x"ec",x"c2",x"87",x"d1"),
  1240 => (x"c2",x"1e",x"7e",x"f8"),
  1241 => (x"eb",x"49",x"d4",x"fa"),
  1242 => (x"86",x"c4",x"87",x"c3"),
  1243 => (x"c5",x"05",x"98",x"70"),
  1244 => (x"c2",x"48",x"c0",x"87"),
  1245 => (x"c0",x"c8",x"87",x"fd"),
  1246 => (x"c4",x"04",x"ad",x"b7"),
  1247 => (x"c4",x"8d",x"4a",x"87"),
  1248 => (x"c0",x"4a",x"75",x"87"),
  1249 => (x"73",x"48",x"6c",x"4d"),
  1250 => (x"58",x"a6",x"c8",x"98"),
  1251 => (x"cc",x"02",x"98",x"70"),
  1252 => (x"73",x"48",x"6c",x"87"),
  1253 => (x"58",x"a6",x"c8",x"98"),
  1254 => (x"f4",x"05",x"98",x"70"),
  1255 => (x"ff",x"7c",x"cd",x"87"),
  1256 => (x"d4",x"c1",x"48",x"d4"),
  1257 => (x"c1",x"49",x"72",x"78"),
  1258 => (x"02",x"99",x"71",x"8a"),
  1259 => (x"97",x"6e",x"87",x"d9"),
  1260 => (x"d4",x"ff",x"48",x"bf"),
  1261 => (x"48",x"6e",x"78",x"08"),
  1262 => (x"a6",x"c4",x"80",x"c1"),
  1263 => (x"c1",x"49",x"72",x"58"),
  1264 => (x"05",x"99",x"71",x"8a"),
  1265 => (x"6c",x"87",x"e7",x"ff"),
  1266 => (x"c4",x"98",x"73",x"48"),
  1267 => (x"98",x"70",x"58",x"a6"),
  1268 => (x"6c",x"87",x"cd",x"02"),
  1269 => (x"c4",x"98",x"73",x"48"),
  1270 => (x"98",x"70",x"58",x"a6"),
  1271 => (x"87",x"f3",x"ff",x"05"),
  1272 => (x"fa",x"c2",x"7c",x"c4"),
  1273 => (x"e1",x"e8",x"49",x"d4"),
  1274 => (x"05",x"9d",x"75",x"87"),
  1275 => (x"6c",x"87",x"ef",x"fd"),
  1276 => (x"c4",x"98",x"73",x"48"),
  1277 => (x"98",x"70",x"58",x"a6"),
  1278 => (x"6c",x"87",x"cd",x"02"),
  1279 => (x"c4",x"98",x"73",x"48"),
  1280 => (x"98",x"70",x"58",x"a6"),
  1281 => (x"87",x"f3",x"ff",x"05"),
  1282 => (x"d4",x"ff",x"7c",x"c5"),
  1283 => (x"78",x"d3",x"c1",x"48"),
  1284 => (x"48",x"6c",x"78",x"c0"),
  1285 => (x"a6",x"c4",x"98",x"73"),
  1286 => (x"02",x"98",x"70",x"58"),
  1287 => (x"48",x"6c",x"87",x"cd"),
  1288 => (x"a6",x"c4",x"98",x"73"),
  1289 => (x"05",x"98",x"70",x"58"),
  1290 => (x"c4",x"87",x"f3",x"ff"),
  1291 => (x"c2",x"48",x"c1",x"7c"),
  1292 => (x"f4",x"48",x"c0",x"87"),
  1293 => (x"87",x"f7",x"f3",x"8e"),
  1294 => (x"6e",x"65",x"70",x"4f"),
  1295 => (x"66",x"20",x"64",x"65"),
  1296 => (x"2c",x"65",x"6c",x"69"),
  1297 => (x"61",x"6f",x"6c",x"20"),
  1298 => (x"67",x"6e",x"69",x"64"),
  1299 => (x"2c",x"73",x"25",x"20"),
  1300 => (x"64",x"69",x"28",x"20"),
  1301 => (x"64",x"25",x"20",x"78"),
  1302 => (x"2e",x"2e",x"2e",x"29"),
  1303 => (x"6f",x"4c",x"00",x"0a"),
  1304 => (x"6e",x"69",x"64",x"61"),
  1305 => (x"2e",x"2e",x"2e",x"67"),
  1306 => (x"6c",x"69",x"46",x"00"),
  1307 => (x"73",x"25",x"20",x"65"),
  1308 => (x"20",x"80",x"00",x"0a"),
  1309 => (x"6b",x"63",x"61",x"42"),
  1310 => (x"61",x"6f",x"4c",x"00"),
  1311 => (x"2e",x"2a",x"20",x"64"),
  1312 => (x"20",x"3a",x"00",x"20"),
  1313 => (x"42",x"20",x"80",x"00"),
  1314 => (x"00",x"6b",x"63",x"61"),
  1315 => (x"78",x"45",x"20",x"80"),
  1316 => (x"49",x"00",x"74",x"69"),
  1317 => (x"69",x"74",x"69",x"6e"),
  1318 => (x"7a",x"69",x"6c",x"61"),
  1319 => (x"20",x"67",x"6e",x"69"),
  1320 => (x"63",x"20",x"44",x"53"),
  1321 => (x"0a",x"64",x"72",x"61"),
  1322 => (x"76",x"61",x"48",x"00"),
  1323 => (x"44",x"53",x"20",x"65"),
  1324 => (x"4f",x"42",x"00",x"0a"),
  1325 => (x"20",x"20",x"54",x"4f"),
  1326 => (x"4f",x"52",x"20",x"20"),
  1327 => (x"5e",x"0e",x"00",x"4d"),
  1328 => (x"0e",x"5d",x"5c",x"5b"),
  1329 => (x"c0",x"4b",x"71",x"1e"),
  1330 => (x"ab",x"b7",x"4d",x"4c"),
  1331 => (x"87",x"e9",x"c0",x"04"),
  1332 => (x"1e",x"e6",x"c5",x"c1"),
  1333 => (x"c4",x"02",x"9d",x"75"),
  1334 => (x"c2",x"4a",x"c0",x"87"),
  1335 => (x"72",x"4a",x"c1",x"87"),
  1336 => (x"87",x"c6",x"e8",x"49"),
  1337 => (x"58",x"a6",x"86",x"c4"),
  1338 => (x"05",x"6e",x"84",x"c1"),
  1339 => (x"4c",x"73",x"87",x"c2"),
  1340 => (x"b7",x"73",x"85",x"c1"),
  1341 => (x"d7",x"ff",x"06",x"ac"),
  1342 => (x"26",x"48",x"6e",x"87"),
  1343 => (x"0e",x"87",x"f0",x"f0"),
  1344 => (x"5d",x"5c",x"5b",x"5e"),
  1345 => (x"4c",x"71",x"1e",x"0e"),
  1346 => (x"e4",x"fa",x"c2",x"49"),
  1347 => (x"ed",x"fe",x"81",x"bf"),
  1348 => (x"1e",x"4d",x"70",x"87"),
  1349 => (x"1e",x"e9",x"d1",x"c1"),
  1350 => (x"87",x"e0",x"ed",x"fe"),
  1351 => (x"9d",x"75",x"86",x"c8"),
  1352 => (x"87",x"fc",x"c0",x"02"),
  1353 => (x"4b",x"c8",x"f5",x"c2"),
  1354 => (x"49",x"cb",x"4a",x"75"),
  1355 => (x"87",x"db",x"f2",x"fe"),
  1356 => (x"91",x"de",x"49",x"74"),
  1357 => (x"48",x"f8",x"fa",x"c2"),
  1358 => (x"a6",x"c4",x"80",x"71"),
  1359 => (x"de",x"d1",x"c1",x"58"),
  1360 => (x"c8",x"49",x"6e",x"48"),
  1361 => (x"41",x"20",x"4a",x"a1"),
  1362 => (x"f9",x"05",x"aa",x"71"),
  1363 => (x"10",x"51",x"10",x"87"),
  1364 => (x"74",x"51",x"10",x"51"),
  1365 => (x"e9",x"c4",x"c1",x"49"),
  1366 => (x"c8",x"f5",x"c2",x"87"),
  1367 => (x"87",x"e3",x"f4",x"49"),
  1368 => (x"49",x"e4",x"f6",x"c1"),
  1369 => (x"87",x"e5",x"c7",x"c1"),
  1370 => (x"87",x"c1",x"c8",x"c1"),
  1371 => (x"87",x"ff",x"ee",x"26"),
  1372 => (x"71",x"1e",x"73",x"1e"),
  1373 => (x"fa",x"c2",x"49",x"4b"),
  1374 => (x"fd",x"81",x"bf",x"e4"),
  1375 => (x"4a",x"70",x"87",x"c0"),
  1376 => (x"87",x"c4",x"02",x"9a"),
  1377 => (x"87",x"df",x"e3",x"49"),
  1378 => (x"48",x"e4",x"fa",x"c2"),
  1379 => (x"49",x"73",x"78",x"c0"),
  1380 => (x"ee",x"87",x"e9",x"c1"),
  1381 => (x"73",x"1e",x"87",x"dd"),
  1382 => (x"c4",x"4b",x"71",x"1e"),
  1383 => (x"c1",x"02",x"4a",x"a3"),
  1384 => (x"8a",x"c1",x"87",x"c8"),
  1385 => (x"8a",x"87",x"dc",x"02"),
  1386 => (x"87",x"f1",x"c0",x"02"),
  1387 => (x"c4",x"c1",x"05",x"8a"),
  1388 => (x"e4",x"fa",x"c2",x"87"),
  1389 => (x"fc",x"c0",x"02",x"bf"),
  1390 => (x"88",x"c1",x"48",x"87"),
  1391 => (x"58",x"e8",x"fa",x"c2"),
  1392 => (x"c2",x"87",x"f2",x"c0"),
  1393 => (x"49",x"bf",x"e4",x"fa"),
  1394 => (x"fa",x"c2",x"89",x"d0"),
  1395 => (x"b7",x"c0",x"59",x"e8"),
  1396 => (x"e0",x"c0",x"03",x"a9"),
  1397 => (x"e4",x"fa",x"c2",x"87"),
  1398 => (x"d8",x"78",x"c0",x"48"),
  1399 => (x"e4",x"fa",x"c2",x"87"),
  1400 => (x"80",x"c1",x"48",x"bf"),
  1401 => (x"58",x"e8",x"fa",x"c2"),
  1402 => (x"fa",x"c2",x"87",x"cb"),
  1403 => (x"d0",x"48",x"bf",x"e4"),
  1404 => (x"e8",x"fa",x"c2",x"80"),
  1405 => (x"c3",x"49",x"73",x"58"),
  1406 => (x"87",x"f7",x"ec",x"87"),
  1407 => (x"5c",x"5b",x"5e",x"0e"),
  1408 => (x"86",x"f0",x"0e",x"5d"),
  1409 => (x"c2",x"59",x"a6",x"d0"),
  1410 => (x"c0",x"4d",x"f8",x"ec"),
  1411 => (x"48",x"a6",x"c4",x"4c"),
  1412 => (x"fa",x"c2",x"78",x"c0"),
  1413 => (x"c0",x"48",x"bf",x"e4"),
  1414 => (x"c1",x"06",x"a8",x"b7"),
  1415 => (x"ec",x"c2",x"87",x"c1"),
  1416 => (x"02",x"98",x"48",x"f8"),
  1417 => (x"c1",x"87",x"f8",x"c0"),
  1418 => (x"c8",x"1e",x"e6",x"c5"),
  1419 => (x"87",x"c7",x"02",x"66"),
  1420 => (x"c0",x"48",x"a6",x"c4"),
  1421 => (x"c4",x"87",x"c5",x"78"),
  1422 => (x"78",x"c1",x"48",x"a6"),
  1423 => (x"e2",x"49",x"66",x"c4"),
  1424 => (x"86",x"c4",x"87",x"e8"),
  1425 => (x"84",x"c1",x"4d",x"70"),
  1426 => (x"c1",x"48",x"66",x"c4"),
  1427 => (x"58",x"a6",x"c8",x"80"),
  1428 => (x"bf",x"e4",x"fa",x"c2"),
  1429 => (x"c6",x"03",x"ac",x"b7"),
  1430 => (x"05",x"9d",x"75",x"87"),
  1431 => (x"c0",x"87",x"c8",x"ff"),
  1432 => (x"02",x"9d",x"75",x"4c"),
  1433 => (x"c1",x"87",x"e3",x"c3"),
  1434 => (x"c8",x"1e",x"e6",x"c5"),
  1435 => (x"87",x"c7",x"02",x"66"),
  1436 => (x"c0",x"48",x"a6",x"cc"),
  1437 => (x"cc",x"87",x"c5",x"78"),
  1438 => (x"78",x"c1",x"48",x"a6"),
  1439 => (x"e1",x"49",x"66",x"cc"),
  1440 => (x"86",x"c4",x"87",x"e8"),
  1441 => (x"02",x"6e",x"58",x"a6"),
  1442 => (x"49",x"87",x"eb",x"c2"),
  1443 => (x"69",x"97",x"81",x"cb"),
  1444 => (x"02",x"99",x"d0",x"49"),
  1445 => (x"c1",x"87",x"d9",x"c1"),
  1446 => (x"74",x"4b",x"f0",x"d5"),
  1447 => (x"c1",x"91",x"cc",x"49"),
  1448 => (x"c8",x"81",x"e4",x"f6"),
  1449 => (x"7a",x"73",x"4a",x"a1"),
  1450 => (x"ff",x"c3",x"81",x"c1"),
  1451 => (x"de",x"49",x"74",x"51"),
  1452 => (x"f8",x"fa",x"c2",x"91"),
  1453 => (x"c2",x"85",x"71",x"4d"),
  1454 => (x"c1",x"7d",x"97",x"c1"),
  1455 => (x"e0",x"c0",x"49",x"a5"),
  1456 => (x"c8",x"f5",x"c2",x"51"),
  1457 => (x"d2",x"02",x"bf",x"97"),
  1458 => (x"c2",x"84",x"c1",x"87"),
  1459 => (x"f5",x"c2",x"4b",x"a5"),
  1460 => (x"49",x"db",x"4a",x"c8"),
  1461 => (x"87",x"f3",x"eb",x"fe"),
  1462 => (x"cd",x"87",x"db",x"c1"),
  1463 => (x"51",x"c0",x"49",x"a5"),
  1464 => (x"a5",x"c2",x"84",x"c1"),
  1465 => (x"cb",x"4a",x"6e",x"4b"),
  1466 => (x"de",x"eb",x"fe",x"49"),
  1467 => (x"87",x"c6",x"c1",x"87"),
  1468 => (x"91",x"cc",x"49",x"74"),
  1469 => (x"81",x"e4",x"f6",x"c1"),
  1470 => (x"d3",x"c1",x"81",x"c8"),
  1471 => (x"f5",x"c2",x"79",x"ff"),
  1472 => (x"02",x"bf",x"97",x"c8"),
  1473 => (x"49",x"74",x"87",x"d8"),
  1474 => (x"84",x"c1",x"91",x"de"),
  1475 => (x"4b",x"f8",x"fa",x"c2"),
  1476 => (x"f5",x"c2",x"83",x"71"),
  1477 => (x"49",x"dd",x"4a",x"c8"),
  1478 => (x"87",x"ef",x"ea",x"fe"),
  1479 => (x"4b",x"74",x"87",x"d8"),
  1480 => (x"fa",x"c2",x"93",x"de"),
  1481 => (x"a3",x"cb",x"83",x"f8"),
  1482 => (x"c1",x"51",x"c0",x"49"),
  1483 => (x"4a",x"6e",x"73",x"84"),
  1484 => (x"ea",x"fe",x"49",x"cb"),
  1485 => (x"66",x"c4",x"87",x"d5"),
  1486 => (x"c8",x"80",x"c1",x"48"),
  1487 => (x"b7",x"c7",x"58",x"a6"),
  1488 => (x"c5",x"c0",x"03",x"ac"),
  1489 => (x"fc",x"05",x"6e",x"87"),
  1490 => (x"b7",x"c7",x"87",x"dd"),
  1491 => (x"d3",x"c0",x"03",x"ac"),
  1492 => (x"de",x"49",x"74",x"87"),
  1493 => (x"f8",x"fa",x"c2",x"91"),
  1494 => (x"c1",x"51",x"c0",x"81"),
  1495 => (x"ac",x"b7",x"c7",x"84"),
  1496 => (x"87",x"ed",x"ff",x"04"),
  1497 => (x"48",x"f9",x"f7",x"c1"),
  1498 => (x"f7",x"c1",x"50",x"c0"),
  1499 => (x"50",x"c2",x"48",x"f8"),
  1500 => (x"48",x"c0",x"f8",x"c1"),
  1501 => (x"78",x"e2",x"de",x"c1"),
  1502 => (x"48",x"fc",x"f7",x"c1"),
  1503 => (x"78",x"f2",x"d1",x"c1"),
  1504 => (x"48",x"cc",x"f8",x"c1"),
  1505 => (x"78",x"d6",x"d6",x"c1"),
  1506 => (x"c0",x"49",x"66",x"cc"),
  1507 => (x"f0",x"87",x"f3",x"fb"),
  1508 => (x"87",x"db",x"e6",x"8e"),
  1509 => (x"c2",x"4a",x"71",x"1e"),
  1510 => (x"72",x"5a",x"d4",x"fa"),
  1511 => (x"87",x"dc",x"f9",x"49"),
  1512 => (x"71",x"1e",x"4f",x"26"),
  1513 => (x"91",x"cc",x"49",x"4a"),
  1514 => (x"81",x"e4",x"f6",x"c1"),
  1515 => (x"48",x"11",x"81",x"c1"),
  1516 => (x"58",x"d0",x"fa",x"c2"),
  1517 => (x"49",x"a2",x"f0",x"c0"),
  1518 => (x"87",x"df",x"e8",x"fe"),
  1519 => (x"dd",x"d5",x"49",x"c0"),
  1520 => (x"0e",x"4f",x"26",x"87"),
  1521 => (x"5d",x"5c",x"5b",x"5e"),
  1522 => (x"71",x"86",x"f0",x"0e"),
  1523 => (x"91",x"cc",x"49",x"4c"),
  1524 => (x"81",x"e4",x"f6",x"c1"),
  1525 => (x"c4",x"7e",x"a1",x"c3"),
  1526 => (x"fa",x"c2",x"48",x"a6"),
  1527 => (x"6e",x"78",x"bf",x"c8"),
  1528 => (x"c4",x"4a",x"bf",x"97"),
  1529 => (x"2b",x"72",x"4b",x"66"),
  1530 => (x"12",x"4a",x"a1",x"c1"),
  1531 => (x"58",x"a6",x"cc",x"48"),
  1532 => (x"83",x"c1",x"9b",x"70"),
  1533 => (x"69",x"97",x"81",x"c2"),
  1534 => (x"04",x"ab",x"b7",x"49"),
  1535 => (x"4b",x"c0",x"87",x"c2"),
  1536 => (x"4a",x"bf",x"97",x"6e"),
  1537 => (x"72",x"49",x"66",x"c8"),
  1538 => (x"c4",x"b9",x"ff",x"31"),
  1539 => (x"4d",x"73",x"99",x"66"),
  1540 => (x"b5",x"71",x"35",x"72"),
  1541 => (x"5d",x"cc",x"fa",x"c2"),
  1542 => (x"c3",x"48",x"d4",x"ff"),
  1543 => (x"d0",x"ff",x"78",x"ff"),
  1544 => (x"c0",x"c8",x"48",x"bf"),
  1545 => (x"a6",x"d0",x"98",x"c0"),
  1546 => (x"02",x"98",x"70",x"58"),
  1547 => (x"d0",x"ff",x"87",x"d0"),
  1548 => (x"c0",x"c8",x"48",x"bf"),
  1549 => (x"a6",x"c4",x"98",x"c0"),
  1550 => (x"05",x"98",x"70",x"58"),
  1551 => (x"d0",x"ff",x"87",x"f0"),
  1552 => (x"78",x"e1",x"c0",x"48"),
  1553 => (x"de",x"48",x"d4",x"ff"),
  1554 => (x"7d",x"0d",x"70",x"78"),
  1555 => (x"c8",x"48",x"75",x"0d"),
  1556 => (x"d4",x"ff",x"28",x"b7"),
  1557 => (x"48",x"75",x"78",x"08"),
  1558 => (x"ff",x"28",x"b7",x"d0"),
  1559 => (x"75",x"78",x"08",x"d4"),
  1560 => (x"28",x"b7",x"d8",x"48"),
  1561 => (x"78",x"08",x"d4",x"ff"),
  1562 => (x"48",x"bf",x"d0",x"ff"),
  1563 => (x"98",x"c0",x"c0",x"c8"),
  1564 => (x"70",x"58",x"a6",x"c4"),
  1565 => (x"87",x"d0",x"02",x"98"),
  1566 => (x"48",x"bf",x"d0",x"ff"),
  1567 => (x"98",x"c0",x"c0",x"c8"),
  1568 => (x"70",x"58",x"a6",x"c4"),
  1569 => (x"87",x"f0",x"05",x"98"),
  1570 => (x"c0",x"48",x"d0",x"ff"),
  1571 => (x"1e",x"c7",x"78",x"e0"),
  1572 => (x"f6",x"c1",x"1e",x"c0"),
  1573 => (x"fa",x"c2",x"1e",x"e4"),
  1574 => (x"c1",x"49",x"bf",x"cc"),
  1575 => (x"49",x"74",x"87",x"e1"),
  1576 => (x"87",x"de",x"f7",x"c0"),
  1577 => (x"c6",x"e2",x"8e",x"e4"),
  1578 => (x"1e",x"73",x"1e",x"87"),
  1579 => (x"fc",x"49",x"4b",x"71"),
  1580 => (x"49",x"73",x"87",x"d1"),
  1581 => (x"e1",x"87",x"cc",x"fc"),
  1582 => (x"73",x"1e",x"87",x"f9"),
  1583 => (x"c2",x"4b",x"71",x"1e"),
  1584 => (x"d5",x"02",x"4a",x"a3"),
  1585 => (x"05",x"8a",x"c1",x"87"),
  1586 => (x"fa",x"c2",x"87",x"db"),
  1587 => (x"d4",x"02",x"bf",x"e0"),
  1588 => (x"88",x"c1",x"48",x"87"),
  1589 => (x"58",x"e4",x"fa",x"c2"),
  1590 => (x"fa",x"c2",x"87",x"cb"),
  1591 => (x"c1",x"48",x"bf",x"e0"),
  1592 => (x"e4",x"fa",x"c2",x"80"),
  1593 => (x"c0",x"1e",x"c7",x"58"),
  1594 => (x"e4",x"f6",x"c1",x"1e"),
  1595 => (x"cc",x"fa",x"c2",x"1e"),
  1596 => (x"87",x"cb",x"49",x"bf"),
  1597 => (x"f6",x"c0",x"49",x"73"),
  1598 => (x"8e",x"f4",x"87",x"c8"),
  1599 => (x"0e",x"87",x"f4",x"e0"),
  1600 => (x"5d",x"5c",x"5b",x"5e"),
  1601 => (x"86",x"d8",x"ff",x"0e"),
  1602 => (x"c8",x"59",x"a6",x"dc"),
  1603 => (x"78",x"c0",x"48",x"a6"),
  1604 => (x"78",x"c0",x"80",x"c4"),
  1605 => (x"c2",x"80",x"c4",x"4d"),
  1606 => (x"78",x"bf",x"e0",x"fa"),
  1607 => (x"c3",x"48",x"d4",x"ff"),
  1608 => (x"d0",x"ff",x"78",x"ff"),
  1609 => (x"c0",x"c8",x"48",x"bf"),
  1610 => (x"a6",x"c4",x"98",x"c0"),
  1611 => (x"02",x"98",x"70",x"58"),
  1612 => (x"d0",x"ff",x"87",x"d0"),
  1613 => (x"c0",x"c8",x"48",x"bf"),
  1614 => (x"a6",x"c4",x"98",x"c0"),
  1615 => (x"05",x"98",x"70",x"58"),
  1616 => (x"d0",x"ff",x"87",x"f0"),
  1617 => (x"78",x"e1",x"c0",x"48"),
  1618 => (x"d4",x"48",x"d4",x"ff"),
  1619 => (x"d5",x"dd",x"ff",x"78"),
  1620 => (x"48",x"d4",x"ff",x"87"),
  1621 => (x"d4",x"78",x"ff",x"c3"),
  1622 => (x"d4",x"ff",x"48",x"a6"),
  1623 => (x"66",x"d4",x"78",x"bf"),
  1624 => (x"a8",x"fb",x"c0",x"48"),
  1625 => (x"87",x"d3",x"c1",x"02"),
  1626 => (x"4a",x"66",x"f8",x"c0"),
  1627 => (x"7e",x"6a",x"82",x"c4"),
  1628 => (x"d1",x"c1",x"1e",x"72"),
  1629 => (x"66",x"c4",x"48",x"f9"),
  1630 => (x"4a",x"a1",x"c8",x"49"),
  1631 => (x"aa",x"71",x"41",x"20"),
  1632 => (x"10",x"87",x"f9",x"05"),
  1633 => (x"c0",x"4a",x"26",x"51"),
  1634 => (x"c8",x"49",x"66",x"f8"),
  1635 => (x"d4",x"de",x"c1",x"81"),
  1636 => (x"c7",x"49",x"6a",x"79"),
  1637 => (x"51",x"66",x"d4",x"81"),
  1638 => (x"1e",x"d8",x"1e",x"c1"),
  1639 => (x"81",x"c8",x"49",x"6a"),
  1640 => (x"87",x"d9",x"dc",x"ff"),
  1641 => (x"66",x"d0",x"86",x"c8"),
  1642 => (x"a8",x"b7",x"c0",x"48"),
  1643 => (x"c1",x"87",x"c4",x"01"),
  1644 => (x"d0",x"87",x"c8",x"4d"),
  1645 => (x"88",x"c1",x"48",x"66"),
  1646 => (x"d4",x"58",x"a6",x"d4"),
  1647 => (x"f4",x"ca",x"02",x"66"),
  1648 => (x"66",x"c0",x"c1",x"87"),
  1649 => (x"ca",x"03",x"ad",x"b7"),
  1650 => (x"d4",x"ff",x"87",x"eb"),
  1651 => (x"78",x"ff",x"c3",x"48"),
  1652 => (x"ff",x"48",x"a6",x"d4"),
  1653 => (x"d4",x"78",x"bf",x"d4"),
  1654 => (x"c6",x"c1",x"48",x"66"),
  1655 => (x"58",x"a6",x"c4",x"88"),
  1656 => (x"c0",x"02",x"98",x"70"),
  1657 => (x"c9",x"48",x"87",x"e6"),
  1658 => (x"58",x"a6",x"c4",x"88"),
  1659 => (x"c4",x"02",x"98",x"70"),
  1660 => (x"c1",x"48",x"87",x"d5"),
  1661 => (x"58",x"a6",x"c4",x"88"),
  1662 => (x"c1",x"02",x"98",x"70"),
  1663 => (x"c4",x"48",x"87",x"e3"),
  1664 => (x"70",x"58",x"a6",x"88"),
  1665 => (x"fe",x"c3",x"02",x"98"),
  1666 => (x"87",x"d3",x"c9",x"87"),
  1667 => (x"c1",x"05",x"66",x"d8"),
  1668 => (x"d4",x"ff",x"87",x"c5"),
  1669 => (x"78",x"ff",x"c3",x"48"),
  1670 => (x"1e",x"ca",x"1e",x"c0"),
  1671 => (x"93",x"cc",x"4b",x"75"),
  1672 => (x"83",x"66",x"c0",x"c1"),
  1673 => (x"6c",x"4c",x"a3",x"c4"),
  1674 => (x"d0",x"da",x"ff",x"49"),
  1675 => (x"de",x"1e",x"c1",x"87"),
  1676 => (x"ff",x"49",x"6c",x"1e"),
  1677 => (x"d0",x"87",x"c6",x"da"),
  1678 => (x"49",x"a3",x"c8",x"86"),
  1679 => (x"79",x"d4",x"de",x"c1"),
  1680 => (x"ad",x"b7",x"66",x"d0"),
  1681 => (x"c1",x"87",x"c5",x"04"),
  1682 => (x"87",x"da",x"c8",x"85"),
  1683 => (x"c1",x"48",x"66",x"d0"),
  1684 => (x"58",x"a6",x"d4",x"88"),
  1685 => (x"ff",x"87",x"cf",x"c8"),
  1686 => (x"d8",x"87",x"cb",x"d9"),
  1687 => (x"c5",x"c8",x"58",x"a6"),
  1688 => (x"d2",x"db",x"ff",x"87"),
  1689 => (x"58",x"a6",x"cc",x"87"),
  1690 => (x"a8",x"b7",x"66",x"cc"),
  1691 => (x"cc",x"87",x"c6",x"06"),
  1692 => (x"66",x"c8",x"48",x"a6"),
  1693 => (x"fe",x"da",x"ff",x"78"),
  1694 => (x"a8",x"ec",x"c0",x"87"),
  1695 => (x"87",x"c7",x"c2",x"05"),
  1696 => (x"c1",x"05",x"66",x"d8"),
  1697 => (x"49",x"75",x"87",x"f7"),
  1698 => (x"f8",x"c0",x"91",x"cc"),
  1699 => (x"a1",x"c4",x"81",x"66"),
  1700 => (x"c1",x"4c",x"6a",x"4a"),
  1701 => (x"66",x"c8",x"4a",x"a1"),
  1702 => (x"79",x"97",x"c2",x"52"),
  1703 => (x"de",x"c1",x"81",x"c8"),
  1704 => (x"d4",x"ff",x"79",x"e2"),
  1705 => (x"78",x"ff",x"c3",x"48"),
  1706 => (x"ff",x"48",x"a6",x"d4"),
  1707 => (x"d4",x"78",x"bf",x"d4"),
  1708 => (x"e8",x"c0",x"02",x"66"),
  1709 => (x"fb",x"c0",x"48",x"87"),
  1710 => (x"e0",x"c0",x"02",x"a8"),
  1711 => (x"97",x"66",x"d4",x"87"),
  1712 => (x"ff",x"84",x"c1",x"7c"),
  1713 => (x"ff",x"c3",x"48",x"d4"),
  1714 => (x"48",x"a6",x"d4",x"78"),
  1715 => (x"78",x"bf",x"d4",x"ff"),
  1716 => (x"c8",x"02",x"66",x"d4"),
  1717 => (x"fb",x"c0",x"48",x"87"),
  1718 => (x"e0",x"ff",x"05",x"a8"),
  1719 => (x"54",x"e0",x"c0",x"87"),
  1720 => (x"c0",x"54",x"c1",x"c2"),
  1721 => (x"66",x"d0",x"7c",x"97"),
  1722 => (x"c5",x"04",x"ad",x"b7"),
  1723 => (x"c5",x"85",x"c1",x"87"),
  1724 => (x"66",x"d0",x"87",x"f4"),
  1725 => (x"d4",x"88",x"c1",x"48"),
  1726 => (x"e9",x"c5",x"58",x"a6"),
  1727 => (x"e5",x"d6",x"ff",x"87"),
  1728 => (x"58",x"a6",x"d8",x"87"),
  1729 => (x"c8",x"87",x"df",x"c5"),
  1730 => (x"66",x"d8",x"48",x"66"),
  1731 => (x"c4",x"c5",x"05",x"a8"),
  1732 => (x"48",x"a6",x"dc",x"87"),
  1733 => (x"d8",x"ff",x"78",x"c0"),
  1734 => (x"a6",x"d8",x"87",x"dd"),
  1735 => (x"d6",x"d8",x"ff",x"58"),
  1736 => (x"a6",x"e4",x"c0",x"87"),
  1737 => (x"a8",x"ec",x"c0",x"58"),
  1738 => (x"87",x"ca",x"c0",x"05"),
  1739 => (x"48",x"a6",x"e0",x"c0"),
  1740 => (x"c0",x"78",x"66",x"d4"),
  1741 => (x"d4",x"ff",x"87",x"c6"),
  1742 => (x"78",x"ff",x"c3",x"48"),
  1743 => (x"91",x"cc",x"49",x"75"),
  1744 => (x"48",x"66",x"f8",x"c0"),
  1745 => (x"a6",x"c4",x"80",x"71"),
  1746 => (x"c3",x"49",x"6e",x"58"),
  1747 => (x"51",x"66",x"d4",x"81"),
  1748 => (x"49",x"66",x"e0",x"c0"),
  1749 => (x"66",x"d4",x"81",x"c1"),
  1750 => (x"71",x"48",x"c1",x"89"),
  1751 => (x"c1",x"49",x"70",x"30"),
  1752 => (x"c1",x"4a",x"6e",x"89"),
  1753 => (x"97",x"09",x"72",x"82"),
  1754 => (x"48",x"6e",x"09",x"79"),
  1755 => (x"fa",x"c2",x"50",x"c2"),
  1756 => (x"d4",x"49",x"bf",x"c8"),
  1757 => (x"97",x"29",x"b7",x"66"),
  1758 => (x"71",x"48",x"4a",x"6a"),
  1759 => (x"a6",x"e8",x"c0",x"98"),
  1760 => (x"c4",x"48",x"6e",x"58"),
  1761 => (x"58",x"a6",x"c8",x"80"),
  1762 => (x"4c",x"bf",x"66",x"c4"),
  1763 => (x"c8",x"48",x"66",x"d8"),
  1764 => (x"c0",x"02",x"a8",x"66"),
  1765 => (x"e0",x"c0",x"87",x"c9"),
  1766 => (x"78",x"c0",x"48",x"a6"),
  1767 => (x"c0",x"87",x"c6",x"c0"),
  1768 => (x"c1",x"48",x"a6",x"e0"),
  1769 => (x"66",x"e0",x"c0",x"78"),
  1770 => (x"1e",x"e0",x"c0",x"1e"),
  1771 => (x"d4",x"ff",x"49",x"74"),
  1772 => (x"86",x"c8",x"87",x"cb"),
  1773 => (x"c0",x"58",x"a6",x"d8"),
  1774 => (x"c1",x"06",x"a8",x"b7"),
  1775 => (x"66",x"d4",x"87",x"da"),
  1776 => (x"bf",x"66",x"c4",x"84"),
  1777 => (x"81",x"e0",x"c0",x"49"),
  1778 => (x"c1",x"4b",x"89",x"74"),
  1779 => (x"71",x"4a",x"c2",x"d2"),
  1780 => (x"87",x"f7",x"d7",x"fe"),
  1781 => (x"66",x"dc",x"84",x"c2"),
  1782 => (x"c0",x"80",x"c1",x"48"),
  1783 => (x"c0",x"58",x"a6",x"e0"),
  1784 => (x"c1",x"49",x"66",x"e4"),
  1785 => (x"02",x"a9",x"70",x"81"),
  1786 => (x"c0",x"87",x"c9",x"c0"),
  1787 => (x"c0",x"48",x"a6",x"e0"),
  1788 => (x"87",x"c6",x"c0",x"78"),
  1789 => (x"48",x"a6",x"e0",x"c0"),
  1790 => (x"e0",x"c0",x"78",x"c1"),
  1791 => (x"66",x"c8",x"1e",x"66"),
  1792 => (x"e0",x"c0",x"49",x"bf"),
  1793 => (x"71",x"89",x"74",x"81"),
  1794 => (x"ff",x"49",x"74",x"1e"),
  1795 => (x"c8",x"87",x"ee",x"d2"),
  1796 => (x"a8",x"b7",x"c0",x"86"),
  1797 => (x"87",x"fe",x"fe",x"01"),
  1798 => (x"c0",x"02",x"66",x"dc"),
  1799 => (x"49",x"6e",x"87",x"d2"),
  1800 => (x"66",x"dc",x"81",x"c2"),
  1801 => (x"c8",x"49",x"6e",x"51"),
  1802 => (x"c3",x"df",x"c1",x"81"),
  1803 => (x"87",x"cd",x"c0",x"79"),
  1804 => (x"81",x"c2",x"49",x"6e"),
  1805 => (x"c8",x"49",x"6e",x"51"),
  1806 => (x"e9",x"e2",x"c1",x"81"),
  1807 => (x"b7",x"66",x"d0",x"79"),
  1808 => (x"c5",x"c0",x"04",x"ad"),
  1809 => (x"c0",x"85",x"c1",x"87"),
  1810 => (x"66",x"d0",x"87",x"dc"),
  1811 => (x"d4",x"88",x"c1",x"48"),
  1812 => (x"d1",x"c0",x"58",x"a6"),
  1813 => (x"cd",x"d1",x"ff",x"87"),
  1814 => (x"58",x"a6",x"d8",x"87"),
  1815 => (x"ff",x"87",x"c7",x"c0"),
  1816 => (x"d8",x"87",x"c3",x"d1"),
  1817 => (x"66",x"d4",x"58",x"a6"),
  1818 => (x"87",x"c9",x"c0",x"02"),
  1819 => (x"b7",x"66",x"c0",x"c1"),
  1820 => (x"d5",x"f5",x"04",x"ad"),
  1821 => (x"ad",x"b7",x"c7",x"87"),
  1822 => (x"87",x"dc",x"c0",x"03"),
  1823 => (x"91",x"cc",x"49",x"75"),
  1824 => (x"81",x"66",x"f8",x"c0"),
  1825 => (x"6a",x"4a",x"a1",x"c4"),
  1826 => (x"c8",x"52",x"c0",x"4a"),
  1827 => (x"c1",x"79",x"c0",x"81"),
  1828 => (x"ad",x"b7",x"c7",x"85"),
  1829 => (x"87",x"e4",x"ff",x"04"),
  1830 => (x"c0",x"02",x"66",x"d8"),
  1831 => (x"f8",x"c0",x"87",x"eb"),
  1832 => (x"d4",x"c1",x"49",x"66"),
  1833 => (x"66",x"f8",x"c0",x"81"),
  1834 => (x"82",x"d5",x"c1",x"4a"),
  1835 => (x"51",x"c2",x"52",x"c0"),
  1836 => (x"49",x"66",x"f8",x"c0"),
  1837 => (x"c1",x"81",x"dc",x"c1"),
  1838 => (x"c0",x"79",x"e2",x"de"),
  1839 => (x"c1",x"49",x"66",x"f8"),
  1840 => (x"d2",x"c1",x"81",x"d8"),
  1841 => (x"d6",x"c0",x"79",x"c5"),
  1842 => (x"66",x"f8",x"c0",x"87"),
  1843 => (x"81",x"d8",x"c1",x"49"),
  1844 => (x"79",x"cc",x"d2",x"c1"),
  1845 => (x"49",x"66",x"f8",x"c0"),
  1846 => (x"c2",x"81",x"dc",x"c1"),
  1847 => (x"c1",x"79",x"ed",x"dd"),
  1848 => (x"c0",x"4a",x"fa",x"e2"),
  1849 => (x"c1",x"49",x"66",x"f8"),
  1850 => (x"79",x"72",x"81",x"e8"),
  1851 => (x"48",x"bf",x"d0",x"ff"),
  1852 => (x"98",x"c0",x"c0",x"c8"),
  1853 => (x"70",x"58",x"a6",x"c4"),
  1854 => (x"d1",x"c0",x"02",x"98"),
  1855 => (x"bf",x"d0",x"ff",x"87"),
  1856 => (x"c0",x"c0",x"c8",x"48"),
  1857 => (x"58",x"a6",x"c4",x"98"),
  1858 => (x"ff",x"05",x"98",x"70"),
  1859 => (x"d0",x"ff",x"87",x"ef"),
  1860 => (x"78",x"e0",x"c0",x"48"),
  1861 => (x"ff",x"48",x"66",x"cc"),
  1862 => (x"d0",x"ff",x"8e",x"d8"),
  1863 => (x"c7",x"1e",x"87",x"d1"),
  1864 => (x"c1",x"1e",x"c0",x"1e"),
  1865 => (x"c2",x"1e",x"e4",x"f6"),
  1866 => (x"49",x"bf",x"cc",x"fa"),
  1867 => (x"c1",x"87",x"d0",x"ef"),
  1868 => (x"c0",x"49",x"e4",x"f6"),
  1869 => (x"f4",x"87",x"d6",x"e8"),
  1870 => (x"1e",x"4f",x"26",x"8e"),
  1871 => (x"c2",x"87",x"c6",x"ca"),
  1872 => (x"c0",x"48",x"e8",x"fa"),
  1873 => (x"48",x"d4",x"ff",x"50"),
  1874 => (x"c1",x"78",x"ff",x"c3"),
  1875 => (x"fe",x"49",x"d3",x"d2"),
  1876 => (x"fe",x"87",x"d4",x"d1"),
  1877 => (x"70",x"87",x"d0",x"de"),
  1878 => (x"87",x"cd",x"02",x"98"),
  1879 => (x"87",x"d0",x"eb",x"fe"),
  1880 => (x"c4",x"02",x"98",x"70"),
  1881 => (x"c2",x"4a",x"c1",x"87"),
  1882 => (x"72",x"4a",x"c0",x"87"),
  1883 => (x"87",x"c8",x"02",x"9a"),
  1884 => (x"49",x"e9",x"d2",x"c1"),
  1885 => (x"87",x"ef",x"d0",x"fe"),
  1886 => (x"bf",x"f8",x"eb",x"c2"),
  1887 => (x"c2",x"d4",x"ff",x"49"),
  1888 => (x"e0",x"fa",x"c2",x"87"),
  1889 => (x"c2",x"78",x"c0",x"48"),
  1890 => (x"c0",x"48",x"cc",x"fa"),
  1891 => (x"cd",x"fe",x"49",x"78"),
  1892 => (x"87",x"dd",x"c3",x"87"),
  1893 => (x"c0",x"87",x"c2",x"c9"),
  1894 => (x"ff",x"87",x"e1",x"e7"),
  1895 => (x"4f",x"26",x"87",x"f6"),
  1896 => (x"00",x"00",x"14",x"b2"),
  1897 => (x"00",x"00",x"00",x"02"),
  1898 => (x"00",x"00",x"2e",x"b8"),
  1899 => (x"00",x"00",x"14",x"ff"),
  1900 => (x"00",x"00",x"00",x"02"),
  1901 => (x"00",x"00",x"2e",x"d6"),
  1902 => (x"00",x"00",x"14",x"ff"),
  1903 => (x"00",x"00",x"00",x"02"),
  1904 => (x"00",x"00",x"2e",x"f4"),
  1905 => (x"00",x"00",x"14",x"ff"),
  1906 => (x"00",x"00",x"00",x"02"),
  1907 => (x"00",x"00",x"2f",x"12"),
  1908 => (x"00",x"00",x"14",x"ff"),
  1909 => (x"00",x"00",x"00",x"02"),
  1910 => (x"00",x"00",x"2f",x"30"),
  1911 => (x"00",x"00",x"14",x"ff"),
  1912 => (x"00",x"00",x"00",x"02"),
  1913 => (x"00",x"00",x"2f",x"4e"),
  1914 => (x"00",x"00",x"14",x"ff"),
  1915 => (x"00",x"00",x"00",x"02"),
  1916 => (x"00",x"00",x"2f",x"6c"),
  1917 => (x"00",x"00",x"14",x"ff"),
  1918 => (x"00",x"00",x"00",x"02"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"00",x"00",x"17",x"a2"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"15",x"96"),
  1924 => (x"d5",x"c1",x"1e",x"1e"),
  1925 => (x"58",x"a6",x"c4",x"87"),
  1926 => (x"1e",x"4f",x"26",x"26"),
  1927 => (x"f0",x"fe",x"4a",x"71"),
  1928 => (x"cd",x"78",x"c0",x"48"),
  1929 => (x"c1",x"0a",x"7a",x"0a"),
  1930 => (x"fe",x"49",x"f1",x"f8"),
  1931 => (x"26",x"87",x"f8",x"cd"),
  1932 => (x"74",x"65",x"53",x"4f"),
  1933 => (x"6e",x"61",x"68",x"20"),
  1934 => (x"72",x"65",x"6c",x"64"),
  1935 => (x"6e",x"49",x"00",x"0a"),
  1936 => (x"74",x"6e",x"69",x"20"),
  1937 => (x"75",x"72",x"72",x"65"),
  1938 => (x"63",x"20",x"74",x"70"),
  1939 => (x"74",x"73",x"6e",x"6f"),
  1940 => (x"74",x"63",x"75",x"72"),
  1941 => (x"00",x"0a",x"72",x"6f"),
  1942 => (x"fe",x"f8",x"c1",x"1e"),
  1943 => (x"c6",x"cd",x"fe",x"49"),
  1944 => (x"d0",x"f8",x"c1",x"87"),
  1945 => (x"87",x"f3",x"fe",x"49"),
  1946 => (x"fe",x"1e",x"4f",x"26"),
  1947 => (x"26",x"48",x"bf",x"f0"),
  1948 => (x"f0",x"fe",x"1e",x"4f"),
  1949 => (x"26",x"78",x"c1",x"48"),
  1950 => (x"f0",x"fe",x"1e",x"4f"),
  1951 => (x"26",x"78",x"c0",x"48"),
  1952 => (x"4a",x"71",x"1e",x"4f"),
  1953 => (x"a2",x"c4",x"7a",x"c0"),
  1954 => (x"c8",x"79",x"c0",x"49"),
  1955 => (x"79",x"c0",x"49",x"a2"),
  1956 => (x"c0",x"49",x"a2",x"cc"),
  1957 => (x"0e",x"4f",x"26",x"79"),
  1958 => (x"0e",x"5c",x"5b",x"5e"),
  1959 => (x"4c",x"71",x"86",x"f8"),
  1960 => (x"cc",x"49",x"a4",x"c8"),
  1961 => (x"48",x"6b",x"4b",x"a4"),
  1962 => (x"a6",x"c4",x"80",x"c1"),
  1963 => (x"c8",x"98",x"cf",x"58"),
  1964 => (x"48",x"69",x"58",x"a6"),
  1965 => (x"05",x"a8",x"66",x"c4"),
  1966 => (x"48",x"6b",x"87",x"d4"),
  1967 => (x"a6",x"c4",x"80",x"c1"),
  1968 => (x"c8",x"98",x"cf",x"58"),
  1969 => (x"48",x"69",x"58",x"a6"),
  1970 => (x"02",x"a8",x"66",x"c4"),
  1971 => (x"e8",x"fe",x"87",x"ec"),
  1972 => (x"a4",x"d0",x"c1",x"87"),
  1973 => (x"c4",x"48",x"6b",x"49"),
  1974 => (x"58",x"a6",x"c4",x"90"),
  1975 => (x"66",x"d4",x"81",x"70"),
  1976 => (x"c1",x"48",x"6b",x"79"),
  1977 => (x"58",x"a6",x"c8",x"80"),
  1978 => (x"7b",x"70",x"98",x"cf"),
  1979 => (x"fd",x"87",x"d2",x"c1"),
  1980 => (x"8e",x"f8",x"87",x"ff"),
  1981 => (x"4d",x"26",x"87",x"c2"),
  1982 => (x"4b",x"26",x"4c",x"26"),
  1983 => (x"5e",x"0e",x"4f",x"26"),
  1984 => (x"0e",x"5d",x"5c",x"5b"),
  1985 => (x"4d",x"71",x"86",x"f8"),
  1986 => (x"6d",x"4c",x"a5",x"c4"),
  1987 => (x"05",x"a8",x"6c",x"48"),
  1988 => (x"48",x"ff",x"87",x"c5"),
  1989 => (x"fd",x"87",x"e5",x"c0"),
  1990 => (x"a5",x"d0",x"87",x"df"),
  1991 => (x"c4",x"48",x"6c",x"4b"),
  1992 => (x"58",x"a6",x"c4",x"90"),
  1993 => (x"4b",x"6b",x"83",x"70"),
  1994 => (x"6c",x"9b",x"ff",x"c3"),
  1995 => (x"c8",x"80",x"c1",x"48"),
  1996 => (x"98",x"cf",x"58",x"a6"),
  1997 => (x"f8",x"fc",x"7c",x"70"),
  1998 => (x"48",x"49",x"73",x"87"),
  1999 => (x"f5",x"fe",x"8e",x"f8"),
  2000 => (x"1e",x"73",x"1e",x"87"),
  2001 => (x"f0",x"fc",x"86",x"f8"),
  2002 => (x"4b",x"bf",x"e0",x"87"),
  2003 => (x"c0",x"e0",x"c0",x"49"),
  2004 => (x"e7",x"c0",x"02",x"99"),
  2005 => (x"c3",x"4a",x"73",x"87"),
  2006 => (x"fe",x"c2",x"9a",x"ff"),
  2007 => (x"c4",x"48",x"bf",x"ca"),
  2008 => (x"58",x"a6",x"c4",x"90"),
  2009 => (x"49",x"da",x"fe",x"c2"),
  2010 => (x"79",x"72",x"81",x"70"),
  2011 => (x"bf",x"ca",x"fe",x"c2"),
  2012 => (x"c8",x"80",x"c1",x"48"),
  2013 => (x"98",x"cf",x"58",x"a6"),
  2014 => (x"58",x"ce",x"fe",x"c2"),
  2015 => (x"c0",x"d0",x"49",x"73"),
  2016 => (x"f2",x"c0",x"02",x"99"),
  2017 => (x"d2",x"fe",x"c2",x"87"),
  2018 => (x"fe",x"c2",x"48",x"bf"),
  2019 => (x"02",x"a8",x"bf",x"d6"),
  2020 => (x"c2",x"87",x"e4",x"c0"),
  2021 => (x"48",x"bf",x"d2",x"fe"),
  2022 => (x"a6",x"c4",x"90",x"c4"),
  2023 => (x"da",x"ff",x"c2",x"58"),
  2024 => (x"e0",x"81",x"70",x"49"),
  2025 => (x"c2",x"78",x"69",x"48"),
  2026 => (x"48",x"bf",x"d2",x"fe"),
  2027 => (x"a6",x"c8",x"80",x"c1"),
  2028 => (x"c2",x"98",x"cf",x"58"),
  2029 => (x"fa",x"58",x"d6",x"fe"),
  2030 => (x"a6",x"c4",x"87",x"f0"),
  2031 => (x"87",x"f1",x"fa",x"58"),
  2032 => (x"f5",x"fc",x"8e",x"f8"),
  2033 => (x"fe",x"c2",x"1e",x"87"),
  2034 => (x"f4",x"fa",x"49",x"ca"),
  2035 => (x"c1",x"fd",x"c1",x"87"),
  2036 => (x"87",x"c7",x"f9",x"49"),
  2037 => (x"26",x"87",x"f5",x"c3"),
  2038 => (x"1e",x"73",x"1e",x"4f"),
  2039 => (x"49",x"ca",x"fe",x"c2"),
  2040 => (x"70",x"87",x"db",x"fc"),
  2041 => (x"aa",x"b7",x"c0",x"4a"),
  2042 => (x"87",x"cc",x"c2",x"04"),
  2043 => (x"05",x"aa",x"f0",x"c3"),
  2044 => (x"c2",x"c2",x"87",x"c9"),
  2045 => (x"78",x"c1",x"48",x"c4"),
  2046 => (x"c3",x"87",x"ed",x"c1"),
  2047 => (x"c9",x"05",x"aa",x"e0"),
  2048 => (x"c8",x"c2",x"c2",x"87"),
  2049 => (x"c1",x"78",x"c1",x"48"),
  2050 => (x"c2",x"c2",x"87",x"de"),
  2051 => (x"c6",x"02",x"bf",x"c8"),
  2052 => (x"a2",x"c0",x"c2",x"87"),
  2053 => (x"72",x"87",x"c2",x"4b"),
  2054 => (x"c4",x"c2",x"c2",x"4b"),
  2055 => (x"e0",x"c0",x"02",x"bf"),
  2056 => (x"c4",x"49",x"73",x"87"),
  2057 => (x"c2",x"91",x"29",x"b7"),
  2058 => (x"73",x"81",x"cc",x"c2"),
  2059 => (x"c2",x"9a",x"cf",x"4a"),
  2060 => (x"72",x"48",x"c1",x"92"),
  2061 => (x"ff",x"4a",x"70",x"30"),
  2062 => (x"69",x"48",x"72",x"ba"),
  2063 => (x"db",x"79",x"70",x"98"),
  2064 => (x"c4",x"49",x"73",x"87"),
  2065 => (x"c2",x"91",x"29",x"b7"),
  2066 => (x"73",x"81",x"cc",x"c2"),
  2067 => (x"c2",x"9a",x"cf",x"4a"),
  2068 => (x"72",x"48",x"c3",x"92"),
  2069 => (x"48",x"4a",x"70",x"30"),
  2070 => (x"79",x"70",x"b0",x"69"),
  2071 => (x"48",x"c8",x"c2",x"c2"),
  2072 => (x"c2",x"c2",x"78",x"c0"),
  2073 => (x"78",x"c0",x"48",x"c4"),
  2074 => (x"49",x"ca",x"fe",x"c2"),
  2075 => (x"70",x"87",x"cf",x"fa"),
  2076 => (x"aa",x"b7",x"c0",x"4a"),
  2077 => (x"87",x"f4",x"fd",x"03"),
  2078 => (x"87",x"c4",x"48",x"c0"),
  2079 => (x"4c",x"26",x"4d",x"26"),
  2080 => (x"4f",x"26",x"4b",x"26"),
  2081 => (x"00",x"00",x"00",x"00"),
  2082 => (x"00",x"00",x"00",x"00"),
  2083 => (x"00",x"00",x"00",x"00"),
  2084 => (x"00",x"00",x"00",x"00"),
  2085 => (x"00",x"00",x"00",x"00"),
  2086 => (x"00",x"00",x"00",x"00"),
  2087 => (x"00",x"00",x"00",x"00"),
  2088 => (x"00",x"00",x"00",x"00"),
  2089 => (x"00",x"00",x"00",x"00"),
  2090 => (x"00",x"00",x"00",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"00",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"00",x"00"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"00",x"00",x"00",x"00"),
  2096 => (x"00",x"00",x"00",x"00"),
  2097 => (x"00",x"00",x"00",x"00"),
  2098 => (x"00",x"00",x"00",x"00"),
  2099 => (x"72",x"4a",x"c0",x"1e"),
  2100 => (x"c2",x"91",x"c4",x"49"),
  2101 => (x"c0",x"81",x"cc",x"c2"),
  2102 => (x"d0",x"82",x"c1",x"79"),
  2103 => (x"ee",x"04",x"aa",x"b7"),
  2104 => (x"0e",x"4f",x"26",x"87"),
  2105 => (x"5d",x"5c",x"5b",x"5e"),
  2106 => (x"f6",x"4d",x"71",x"0e"),
  2107 => (x"4a",x"75",x"87",x"cb"),
  2108 => (x"92",x"2a",x"b7",x"c4"),
  2109 => (x"82",x"cc",x"c2",x"c2"),
  2110 => (x"9c",x"cf",x"4c",x"75"),
  2111 => (x"49",x"6a",x"94",x"c2"),
  2112 => (x"c3",x"2b",x"74",x"4b"),
  2113 => (x"74",x"48",x"c2",x"9b"),
  2114 => (x"ff",x"4c",x"70",x"30"),
  2115 => (x"71",x"48",x"74",x"bc"),
  2116 => (x"f5",x"7a",x"70",x"98"),
  2117 => (x"48",x"73",x"87",x"db"),
  2118 => (x"1e",x"87",x"e1",x"fd"),
  2119 => (x"bf",x"d0",x"ff",x"1e"),
  2120 => (x"c0",x"c0",x"c8",x"48"),
  2121 => (x"58",x"a6",x"c4",x"98"),
  2122 => (x"d0",x"02",x"98",x"70"),
  2123 => (x"bf",x"d0",x"ff",x"87"),
  2124 => (x"c0",x"c0",x"c8",x"48"),
  2125 => (x"58",x"a6",x"c4",x"98"),
  2126 => (x"f0",x"05",x"98",x"70"),
  2127 => (x"48",x"d0",x"ff",x"87"),
  2128 => (x"71",x"78",x"e1",x"c4"),
  2129 => (x"08",x"d4",x"ff",x"48"),
  2130 => (x"48",x"66",x"c8",x"78"),
  2131 => (x"78",x"08",x"d4",x"ff"),
  2132 => (x"1e",x"4f",x"26",x"26"),
  2133 => (x"c8",x"4a",x"71",x"1e"),
  2134 => (x"72",x"1e",x"49",x"66"),
  2135 => (x"87",x"fb",x"fe",x"49"),
  2136 => (x"d0",x"ff",x"86",x"c4"),
  2137 => (x"c0",x"c8",x"48",x"bf"),
  2138 => (x"a6",x"c4",x"98",x"c0"),
  2139 => (x"02",x"98",x"70",x"58"),
  2140 => (x"d0",x"ff",x"87",x"d0"),
  2141 => (x"c0",x"c8",x"48",x"bf"),
  2142 => (x"a6",x"c4",x"98",x"c0"),
  2143 => (x"05",x"98",x"70",x"58"),
  2144 => (x"d0",x"ff",x"87",x"f0"),
  2145 => (x"78",x"e0",x"c0",x"48"),
  2146 => (x"1e",x"4f",x"26",x"26"),
  2147 => (x"4b",x"71",x"1e",x"73"),
  2148 => (x"73",x"1e",x"66",x"c8"),
  2149 => (x"a2",x"e0",x"c1",x"4a"),
  2150 => (x"87",x"f7",x"fe",x"49"),
  2151 => (x"26",x"87",x"c4",x"26"),
  2152 => (x"26",x"4c",x"26",x"4d"),
  2153 => (x"1e",x"4f",x"26",x"4b"),
  2154 => (x"bf",x"d0",x"ff",x"1e"),
  2155 => (x"c0",x"c0",x"c8",x"48"),
  2156 => (x"58",x"a6",x"c4",x"98"),
  2157 => (x"d0",x"02",x"98",x"70"),
  2158 => (x"bf",x"d0",x"ff",x"87"),
  2159 => (x"c0",x"c0",x"c8",x"48"),
  2160 => (x"58",x"a6",x"c4",x"98"),
  2161 => (x"f0",x"05",x"98",x"70"),
  2162 => (x"48",x"d0",x"ff",x"87"),
  2163 => (x"71",x"78",x"c9",x"c4"),
  2164 => (x"08",x"d4",x"ff",x"48"),
  2165 => (x"4f",x"26",x"26",x"78"),
  2166 => (x"4a",x"71",x"1e",x"1e"),
  2167 => (x"87",x"c7",x"ff",x"49"),
  2168 => (x"48",x"bf",x"d0",x"ff"),
  2169 => (x"98",x"c0",x"c0",x"c8"),
  2170 => (x"70",x"58",x"a6",x"c4"),
  2171 => (x"87",x"d0",x"02",x"98"),
  2172 => (x"48",x"bf",x"d0",x"ff"),
  2173 => (x"98",x"c0",x"c0",x"c8"),
  2174 => (x"70",x"58",x"a6",x"c4"),
  2175 => (x"87",x"f0",x"05",x"98"),
  2176 => (x"c8",x"48",x"d0",x"ff"),
  2177 => (x"4f",x"26",x"26",x"78"),
  2178 => (x"1e",x"1e",x"73",x"1e"),
  2179 => (x"c0",x"c3",x"4b",x"71"),
  2180 => (x"c3",x"02",x"bf",x"e6"),
  2181 => (x"87",x"cc",x"c3",x"87"),
  2182 => (x"48",x"bf",x"d0",x"ff"),
  2183 => (x"98",x"c0",x"c0",x"c8"),
  2184 => (x"70",x"58",x"a6",x"c4"),
  2185 => (x"87",x"d0",x"02",x"98"),
  2186 => (x"48",x"bf",x"d0",x"ff"),
  2187 => (x"98",x"c0",x"c0",x"c8"),
  2188 => (x"70",x"58",x"a6",x"c4"),
  2189 => (x"87",x"f0",x"05",x"98"),
  2190 => (x"c4",x"48",x"d0",x"ff"),
  2191 => (x"48",x"73",x"78",x"c9"),
  2192 => (x"ff",x"b0",x"e0",x"c0"),
  2193 => (x"c3",x"78",x"08",x"d4"),
  2194 => (x"c0",x"48",x"da",x"c0"),
  2195 => (x"02",x"66",x"cc",x"78"),
  2196 => (x"ff",x"c3",x"87",x"c5"),
  2197 => (x"c0",x"87",x"c2",x"49"),
  2198 => (x"e2",x"c0",x"c3",x"49"),
  2199 => (x"02",x"66",x"d0",x"59"),
  2200 => (x"d5",x"c5",x"87",x"c6"),
  2201 => (x"87",x"c4",x"4a",x"d5"),
  2202 => (x"4a",x"ff",x"ff",x"cf"),
  2203 => (x"5a",x"e6",x"c0",x"c3"),
  2204 => (x"48",x"e6",x"c0",x"c3"),
  2205 => (x"c4",x"26",x"78",x"c1"),
  2206 => (x"26",x"4d",x"26",x"87"),
  2207 => (x"26",x"4b",x"26",x"4c"),
  2208 => (x"5b",x"5e",x"0e",x"4f"),
  2209 => (x"71",x"0e",x"5d",x"5c"),
  2210 => (x"e2",x"c0",x"c3",x"4a"),
  2211 => (x"9a",x"72",x"4c",x"bf"),
  2212 => (x"49",x"87",x"cb",x"02"),
  2213 => (x"c9",x"c2",x"91",x"c8"),
  2214 => (x"83",x"71",x"4b",x"c2"),
  2215 => (x"cd",x"c2",x"87",x"c4"),
  2216 => (x"4d",x"c0",x"4b",x"c2"),
  2217 => (x"99",x"74",x"49",x"13"),
  2218 => (x"bf",x"de",x"c0",x"c3"),
  2219 => (x"ff",x"b8",x"71",x"48"),
  2220 => (x"c1",x"78",x"08",x"d4"),
  2221 => (x"c8",x"85",x"2c",x"b7"),
  2222 => (x"e7",x"04",x"ad",x"b7"),
  2223 => (x"da",x"c0",x"c3",x"87"),
  2224 => (x"80",x"c8",x"48",x"bf"),
  2225 => (x"58",x"de",x"c0",x"c3"),
  2226 => (x"1e",x"87",x"ee",x"fe"),
  2227 => (x"4b",x"71",x"1e",x"73"),
  2228 => (x"02",x"9a",x"4a",x"13"),
  2229 => (x"49",x"72",x"87",x"cb"),
  2230 => (x"13",x"87",x"e6",x"fe"),
  2231 => (x"f5",x"05",x"9a",x"4a"),
  2232 => (x"87",x"d9",x"fe",x"87"),
  2233 => (x"c0",x"c3",x"1e",x"1e"),
  2234 => (x"c3",x"49",x"bf",x"da"),
  2235 => (x"c1",x"48",x"da",x"c0"),
  2236 => (x"c0",x"c4",x"78",x"a1"),
  2237 => (x"db",x"03",x"a9",x"b7"),
  2238 => (x"48",x"d4",x"ff",x"87"),
  2239 => (x"bf",x"de",x"c0",x"c3"),
  2240 => (x"da",x"c0",x"c3",x"78"),
  2241 => (x"c0",x"c3",x"49",x"bf"),
  2242 => (x"a1",x"c1",x"48",x"da"),
  2243 => (x"b7",x"c0",x"c4",x"78"),
  2244 => (x"87",x"e5",x"04",x"a9"),
  2245 => (x"48",x"bf",x"d0",x"ff"),
  2246 => (x"98",x"c0",x"c0",x"c8"),
  2247 => (x"70",x"58",x"a6",x"c4"),
  2248 => (x"87",x"d0",x"02",x"98"),
  2249 => (x"48",x"bf",x"d0",x"ff"),
  2250 => (x"98",x"c0",x"c0",x"c8"),
  2251 => (x"70",x"58",x"a6",x"c4"),
  2252 => (x"87",x"f0",x"05",x"98"),
  2253 => (x"c8",x"48",x"d0",x"ff"),
  2254 => (x"e6",x"c0",x"c3",x"78"),
  2255 => (x"26",x"78",x"c0",x"48"),
  2256 => (x"00",x"00",x"4f",x"26"),
  2257 => (x"00",x"00",x"00",x"00"),
  2258 => (x"00",x"00",x"00",x"00"),
  2259 => (x"00",x"5f",x"5f",x"00"),
  2260 => (x"03",x"00",x"00",x"00"),
  2261 => (x"03",x"03",x"00",x"03"),
  2262 => (x"7f",x"14",x"00",x"00"),
  2263 => (x"7f",x"7f",x"14",x"7f"),
  2264 => (x"24",x"00",x"00",x"14"),
  2265 => (x"3a",x"6b",x"6b",x"2e"),
  2266 => (x"6a",x"4c",x"00",x"12"),
  2267 => (x"56",x"6c",x"18",x"36"),
  2268 => (x"7e",x"30",x"00",x"32"),
  2269 => (x"3a",x"77",x"59",x"4f"),
  2270 => (x"00",x"00",x"40",x"68"),
  2271 => (x"00",x"03",x"07",x"04"),
  2272 => (x"00",x"00",x"00",x"00"),
  2273 => (x"41",x"63",x"3e",x"1c"),
  2274 => (x"00",x"00",x"00",x"00"),
  2275 => (x"1c",x"3e",x"63",x"41"),
  2276 => (x"2a",x"08",x"00",x"00"),
  2277 => (x"3e",x"1c",x"1c",x"3e"),
  2278 => (x"08",x"00",x"08",x"2a"),
  2279 => (x"08",x"3e",x"3e",x"08"),
  2280 => (x"00",x"00",x"00",x"08"),
  2281 => (x"00",x"60",x"e0",x"80"),
  2282 => (x"08",x"00",x"00",x"00"),
  2283 => (x"08",x"08",x"08",x"08"),
  2284 => (x"00",x"00",x"00",x"08"),
  2285 => (x"00",x"60",x"60",x"00"),
  2286 => (x"60",x"40",x"00",x"00"),
  2287 => (x"06",x"0c",x"18",x"30"),
  2288 => (x"3e",x"00",x"01",x"03"),
  2289 => (x"7f",x"4d",x"59",x"7f"),
  2290 => (x"04",x"00",x"00",x"3e"),
  2291 => (x"00",x"7f",x"7f",x"06"),
  2292 => (x"42",x"00",x"00",x"00"),
  2293 => (x"4f",x"59",x"71",x"63"),
  2294 => (x"22",x"00",x"00",x"46"),
  2295 => (x"7f",x"49",x"49",x"63"),
  2296 => (x"1c",x"18",x"00",x"36"),
  2297 => (x"7f",x"7f",x"13",x"16"),
  2298 => (x"27",x"00",x"00",x"10"),
  2299 => (x"7d",x"45",x"45",x"67"),
  2300 => (x"3c",x"00",x"00",x"39"),
  2301 => (x"79",x"49",x"4b",x"7e"),
  2302 => (x"01",x"00",x"00",x"30"),
  2303 => (x"0f",x"79",x"71",x"01"),
  2304 => (x"36",x"00",x"00",x"07"),
  2305 => (x"7f",x"49",x"49",x"7f"),
  2306 => (x"06",x"00",x"00",x"36"),
  2307 => (x"3f",x"69",x"49",x"4f"),
  2308 => (x"00",x"00",x"00",x"1e"),
  2309 => (x"00",x"66",x"66",x"00"),
  2310 => (x"00",x"00",x"00",x"00"),
  2311 => (x"00",x"66",x"e6",x"80"),
  2312 => (x"08",x"00",x"00",x"00"),
  2313 => (x"22",x"14",x"14",x"08"),
  2314 => (x"14",x"00",x"00",x"22"),
  2315 => (x"14",x"14",x"14",x"14"),
  2316 => (x"22",x"00",x"00",x"14"),
  2317 => (x"08",x"14",x"14",x"22"),
  2318 => (x"02",x"00",x"00",x"08"),
  2319 => (x"0f",x"59",x"51",x"03"),
  2320 => (x"7f",x"3e",x"00",x"06"),
  2321 => (x"1f",x"55",x"5d",x"41"),
  2322 => (x"7e",x"00",x"00",x"1e"),
  2323 => (x"7f",x"09",x"09",x"7f"),
  2324 => (x"7f",x"00",x"00",x"7e"),
  2325 => (x"7f",x"49",x"49",x"7f"),
  2326 => (x"1c",x"00",x"00",x"36"),
  2327 => (x"41",x"41",x"63",x"3e"),
  2328 => (x"7f",x"00",x"00",x"41"),
  2329 => (x"3e",x"63",x"41",x"7f"),
  2330 => (x"7f",x"00",x"00",x"1c"),
  2331 => (x"41",x"49",x"49",x"7f"),
  2332 => (x"7f",x"00",x"00",x"41"),
  2333 => (x"01",x"09",x"09",x"7f"),
  2334 => (x"3e",x"00",x"00",x"01"),
  2335 => (x"7b",x"49",x"41",x"7f"),
  2336 => (x"7f",x"00",x"00",x"7a"),
  2337 => (x"7f",x"08",x"08",x"7f"),
  2338 => (x"00",x"00",x"00",x"7f"),
  2339 => (x"41",x"7f",x"7f",x"41"),
  2340 => (x"20",x"00",x"00",x"00"),
  2341 => (x"7f",x"40",x"40",x"60"),
  2342 => (x"7f",x"7f",x"00",x"3f"),
  2343 => (x"63",x"36",x"1c",x"08"),
  2344 => (x"7f",x"00",x"00",x"41"),
  2345 => (x"40",x"40",x"40",x"7f"),
  2346 => (x"7f",x"7f",x"00",x"40"),
  2347 => (x"7f",x"06",x"0c",x"06"),
  2348 => (x"7f",x"7f",x"00",x"7f"),
  2349 => (x"7f",x"18",x"0c",x"06"),
  2350 => (x"3e",x"00",x"00",x"7f"),
  2351 => (x"7f",x"41",x"41",x"7f"),
  2352 => (x"7f",x"00",x"00",x"3e"),
  2353 => (x"0f",x"09",x"09",x"7f"),
  2354 => (x"7f",x"3e",x"00",x"06"),
  2355 => (x"7e",x"7f",x"61",x"41"),
  2356 => (x"7f",x"00",x"00",x"40"),
  2357 => (x"7f",x"19",x"09",x"7f"),
  2358 => (x"26",x"00",x"00",x"66"),
  2359 => (x"7b",x"59",x"4d",x"6f"),
  2360 => (x"01",x"00",x"00",x"32"),
  2361 => (x"01",x"7f",x"7f",x"01"),
  2362 => (x"3f",x"00",x"00",x"01"),
  2363 => (x"7f",x"40",x"40",x"7f"),
  2364 => (x"0f",x"00",x"00",x"3f"),
  2365 => (x"3f",x"70",x"70",x"3f"),
  2366 => (x"7f",x"7f",x"00",x"0f"),
  2367 => (x"7f",x"30",x"18",x"30"),
  2368 => (x"63",x"41",x"00",x"7f"),
  2369 => (x"36",x"1c",x"1c",x"36"),
  2370 => (x"03",x"01",x"41",x"63"),
  2371 => (x"06",x"7c",x"7c",x"06"),
  2372 => (x"71",x"61",x"01",x"03"),
  2373 => (x"43",x"47",x"4d",x"59"),
  2374 => (x"00",x"00",x"00",x"41"),
  2375 => (x"41",x"41",x"7f",x"7f"),
  2376 => (x"03",x"01",x"00",x"00"),
  2377 => (x"30",x"18",x"0c",x"06"),
  2378 => (x"00",x"00",x"40",x"60"),
  2379 => (x"7f",x"7f",x"41",x"41"),
  2380 => (x"0c",x"08",x"00",x"00"),
  2381 => (x"0c",x"06",x"03",x"06"),
  2382 => (x"80",x"80",x"00",x"08"),
  2383 => (x"80",x"80",x"80",x"80"),
  2384 => (x"00",x"00",x"00",x"80"),
  2385 => (x"04",x"07",x"03",x"00"),
  2386 => (x"20",x"00",x"00",x"00"),
  2387 => (x"7c",x"54",x"54",x"74"),
  2388 => (x"7f",x"00",x"00",x"78"),
  2389 => (x"7c",x"44",x"44",x"7f"),
  2390 => (x"38",x"00",x"00",x"38"),
  2391 => (x"44",x"44",x"44",x"7c"),
  2392 => (x"38",x"00",x"00",x"00"),
  2393 => (x"7f",x"44",x"44",x"7c"),
  2394 => (x"38",x"00",x"00",x"7f"),
  2395 => (x"5c",x"54",x"54",x"7c"),
  2396 => (x"04",x"00",x"00",x"18"),
  2397 => (x"05",x"05",x"7f",x"7e"),
  2398 => (x"18",x"00",x"00",x"00"),
  2399 => (x"fc",x"a4",x"a4",x"bc"),
  2400 => (x"7f",x"00",x"00",x"7c"),
  2401 => (x"7c",x"04",x"04",x"7f"),
  2402 => (x"00",x"00",x"00",x"78"),
  2403 => (x"40",x"7d",x"3d",x"00"),
  2404 => (x"80",x"00",x"00",x"00"),
  2405 => (x"7d",x"fd",x"80",x"80"),
  2406 => (x"7f",x"00",x"00",x"00"),
  2407 => (x"6c",x"38",x"10",x"7f"),
  2408 => (x"00",x"00",x"00",x"44"),
  2409 => (x"40",x"7f",x"3f",x"00"),
  2410 => (x"7c",x"7c",x"00",x"00"),
  2411 => (x"7c",x"0c",x"18",x"0c"),
  2412 => (x"7c",x"00",x"00",x"78"),
  2413 => (x"7c",x"04",x"04",x"7c"),
  2414 => (x"38",x"00",x"00",x"78"),
  2415 => (x"7c",x"44",x"44",x"7c"),
  2416 => (x"fc",x"00",x"00",x"38"),
  2417 => (x"3c",x"24",x"24",x"fc"),
  2418 => (x"18",x"00",x"00",x"18"),
  2419 => (x"fc",x"24",x"24",x"3c"),
  2420 => (x"7c",x"00",x"00",x"fc"),
  2421 => (x"0c",x"04",x"04",x"7c"),
  2422 => (x"48",x"00",x"00",x"08"),
  2423 => (x"74",x"54",x"54",x"5c"),
  2424 => (x"04",x"00",x"00",x"20"),
  2425 => (x"44",x"44",x"7f",x"3f"),
  2426 => (x"3c",x"00",x"00",x"00"),
  2427 => (x"7c",x"40",x"40",x"7c"),
  2428 => (x"1c",x"00",x"00",x"7c"),
  2429 => (x"3c",x"60",x"60",x"3c"),
  2430 => (x"7c",x"3c",x"00",x"1c"),
  2431 => (x"7c",x"60",x"30",x"60"),
  2432 => (x"6c",x"44",x"00",x"3c"),
  2433 => (x"6c",x"38",x"10",x"38"),
  2434 => (x"1c",x"00",x"00",x"44"),
  2435 => (x"3c",x"60",x"e0",x"bc"),
  2436 => (x"44",x"00",x"00",x"1c"),
  2437 => (x"4c",x"5c",x"74",x"64"),
  2438 => (x"08",x"00",x"00",x"44"),
  2439 => (x"41",x"77",x"3e",x"08"),
  2440 => (x"00",x"00",x"00",x"41"),
  2441 => (x"00",x"7f",x"7f",x"00"),
  2442 => (x"41",x"00",x"00",x"00"),
  2443 => (x"08",x"3e",x"77",x"41"),
  2444 => (x"01",x"02",x"00",x"08"),
  2445 => (x"02",x"02",x"03",x"01"),
  2446 => (x"7f",x"7f",x"00",x"01"),
  2447 => (x"7f",x"7f",x"7f",x"7f"),
  2448 => (x"08",x"08",x"00",x"7f"),
  2449 => (x"3e",x"3e",x"1c",x"1c"),
  2450 => (x"7f",x"7f",x"7f",x"7f"),
  2451 => (x"1c",x"1c",x"3e",x"3e"),
  2452 => (x"10",x"00",x"08",x"08"),
  2453 => (x"18",x"7c",x"7c",x"18"),
  2454 => (x"10",x"00",x"00",x"10"),
  2455 => (x"30",x"7c",x"7c",x"30"),
  2456 => (x"30",x"10",x"00",x"10"),
  2457 => (x"1e",x"78",x"60",x"60"),
  2458 => (x"66",x"42",x"00",x"06"),
  2459 => (x"66",x"3c",x"18",x"3c"),
  2460 => (x"38",x"78",x"00",x"42"),
  2461 => (x"6c",x"c6",x"c2",x"6a"),
  2462 => (x"00",x"60",x"00",x"38"),
  2463 => (x"00",x"00",x"60",x"00"),
  2464 => (x"5e",x"0e",x"00",x"60"),
  2465 => (x"0e",x"5d",x"5c",x"5b"),
  2466 => (x"c3",x"4c",x"71",x"1e"),
  2467 => (x"4b",x"bf",x"ee",x"c0"),
  2468 => (x"48",x"f2",x"c0",x"c3"),
  2469 => (x"1e",x"74",x"78",x"c0"),
  2470 => (x"1e",x"dd",x"dc",x"c2"),
  2471 => (x"87",x"dc",x"e7",x"fd"),
  2472 => (x"6b",x"97",x"86",x"c8"),
  2473 => (x"c1",x"02",x"99",x"49"),
  2474 => (x"1e",x"c0",x"87",x"c6"),
  2475 => (x"c3",x"48",x"a6",x"c4"),
  2476 => (x"78",x"bf",x"f2",x"c0"),
  2477 => (x"02",x"ac",x"66",x"c4"),
  2478 => (x"4d",x"c0",x"87",x"c4"),
  2479 => (x"4d",x"c1",x"87",x"c2"),
  2480 => (x"66",x"c8",x"1e",x"75"),
  2481 => (x"87",x"c0",x"ed",x"49"),
  2482 => (x"e0",x"c0",x"86",x"c8"),
  2483 => (x"87",x"f1",x"ee",x"49"),
  2484 => (x"6a",x"4a",x"a3",x"c4"),
  2485 => (x"87",x"f3",x"ef",x"49"),
  2486 => (x"c3",x"87",x"c9",x"f0"),
  2487 => (x"48",x"bf",x"f2",x"c0"),
  2488 => (x"c0",x"c3",x"80",x"c1"),
  2489 => (x"83",x"cc",x"58",x"f6"),
  2490 => (x"99",x"49",x"6b",x"97"),
  2491 => (x"87",x"fa",x"fe",x"05"),
  2492 => (x"bf",x"f2",x"c0",x"c3"),
  2493 => (x"ad",x"b7",x"c8",x"4d"),
  2494 => (x"c0",x"87",x"d9",x"03"),
  2495 => (x"c0",x"c3",x"1e",x"1e"),
  2496 => (x"ec",x"49",x"bf",x"f2"),
  2497 => (x"86",x"c8",x"87",x"c2"),
  2498 => (x"c1",x"87",x"d9",x"ef"),
  2499 => (x"ad",x"b7",x"c8",x"85"),
  2500 => (x"87",x"e7",x"ff",x"04"),
  2501 => (x"26",x"4d",x"26",x"26"),
  2502 => (x"26",x"4b",x"26",x"4c"),
  2503 => (x"67",x"69",x"48",x"4f"),
  2504 => (x"67",x"69",x"6c",x"68"),
  2505 => (x"72",x"20",x"74",x"68"),
  2506 => (x"25",x"20",x"77",x"6f"),
  2507 => (x"4d",x"00",x"0a",x"64"),
  2508 => (x"20",x"75",x"6e",x"65"),
  2509 => (x"69",x"73",x"69",x"76"),
  2510 => (x"20",x"65",x"6c",x"62"),
  2511 => (x"00",x"0a",x"64",x"25"),
  2512 => (x"6c",x"6c",x"61",x"43"),
  2513 => (x"6b",x"63",x"61",x"62"),
  2514 => (x"0a",x"78",x"25",x"20"),
  2515 => (x"4a",x"71",x"1e",x"00"),
  2516 => (x"5a",x"f2",x"c0",x"c3"),
  2517 => (x"bf",x"f6",x"c0",x"c3"),
  2518 => (x"87",x"e6",x"fc",x"49"),
  2519 => (x"bf",x"f2",x"c0",x"c3"),
  2520 => (x"c3",x"89",x"c1",x"49"),
  2521 => (x"71",x"59",x"fa",x"c0"),
  2522 => (x"26",x"87",x"d7",x"fc"),
  2523 => (x"c0",x"c1",x"1e",x"4f"),
  2524 => (x"87",x"e4",x"e9",x"49"),
  2525 => (x"48",x"e1",x"eb",x"c2"),
  2526 => (x"4f",x"26",x"78",x"c0"),
  2527 => (x"5c",x"5b",x"5e",x"0e"),
  2528 => (x"86",x"f4",x"0e",x"5d"),
  2529 => (x"c0",x"48",x"a6",x"c8"),
  2530 => (x"7e",x"bf",x"ec",x"78"),
  2531 => (x"c0",x"c3",x"80",x"fc"),
  2532 => (x"c3",x"78",x"bf",x"ee"),
  2533 => (x"4d",x"bf",x"fa",x"c0"),
  2534 => (x"c7",x"4c",x"bf",x"e8"),
  2535 => (x"87",x"c3",x"e5",x"49"),
  2536 => (x"99",x"c2",x"49",x"70"),
  2537 => (x"c2",x"87",x"cf",x"05"),
  2538 => (x"49",x"bf",x"d9",x"eb"),
  2539 => (x"99",x"6e",x"b9",x"ff"),
  2540 => (x"c0",x"02",x"99",x"c1"),
  2541 => (x"49",x"c7",x"87",x"fd"),
  2542 => (x"70",x"87",x"e8",x"e4"),
  2543 => (x"87",x"cd",x"02",x"98"),
  2544 => (x"c7",x"87",x"d6",x"e0"),
  2545 => (x"87",x"db",x"e4",x"49"),
  2546 => (x"f3",x"05",x"98",x"70"),
  2547 => (x"e1",x"eb",x"c2",x"87"),
  2548 => (x"dc",x"c2",x"1e",x"bf"),
  2549 => (x"e2",x"fd",x"1e",x"ef"),
  2550 => (x"86",x"c8",x"87",x"e2"),
  2551 => (x"bf",x"e1",x"eb",x"c2"),
  2552 => (x"c2",x"ba",x"c1",x"4a"),
  2553 => (x"c1",x"5a",x"e5",x"eb"),
  2554 => (x"e7",x"49",x"a2",x"c0"),
  2555 => (x"a6",x"c8",x"87",x"ea"),
  2556 => (x"c2",x"78",x"c1",x"48"),
  2557 => (x"6e",x"48",x"d9",x"eb"),
  2558 => (x"e1",x"eb",x"c2",x"78"),
  2559 => (x"da",x"c1",x"05",x"bf"),
  2560 => (x"48",x"a6",x"c4",x"87"),
  2561 => (x"78",x"c0",x"c0",x"c8"),
  2562 => (x"7e",x"e5",x"eb",x"c2"),
  2563 => (x"49",x"bf",x"97",x"6e"),
  2564 => (x"80",x"c1",x"48",x"6e"),
  2565 => (x"71",x"58",x"a6",x"c4"),
  2566 => (x"70",x"87",x"c8",x"e3"),
  2567 => (x"87",x"c3",x"02",x"98"),
  2568 => (x"c4",x"b4",x"66",x"c4"),
  2569 => (x"b7",x"c1",x"48",x"66"),
  2570 => (x"58",x"a6",x"c8",x"28"),
  2571 => (x"ff",x"05",x"98",x"70"),
  2572 => (x"49",x"74",x"87",x"da"),
  2573 => (x"71",x"99",x"ff",x"c3"),
  2574 => (x"e5",x"49",x"c0",x"1e"),
  2575 => (x"49",x"74",x"87",x"cd"),
  2576 => (x"71",x"29",x"b7",x"c8"),
  2577 => (x"e5",x"49",x"c1",x"1e"),
  2578 => (x"86",x"c8",x"87",x"c1"),
  2579 => (x"e2",x"49",x"fd",x"c3"),
  2580 => (x"fa",x"c3",x"87",x"d1"),
  2581 => (x"87",x"cb",x"e2",x"49"),
  2582 => (x"74",x"87",x"e9",x"c9"),
  2583 => (x"99",x"ff",x"c3",x"49"),
  2584 => (x"71",x"2c",x"b7",x"c8"),
  2585 => (x"02",x"9c",x"74",x"b4"),
  2586 => (x"c8",x"ff",x"87",x"df"),
  2587 => (x"49",x"6e",x"7e",x"bf"),
  2588 => (x"bf",x"dd",x"eb",x"c2"),
  2589 => (x"a9",x"c0",x"c2",x"89"),
  2590 => (x"87",x"c4",x"c0",x"03"),
  2591 => (x"87",x"cf",x"4c",x"c0"),
  2592 => (x"48",x"dd",x"eb",x"c2"),
  2593 => (x"c6",x"c0",x"78",x"6e"),
  2594 => (x"dd",x"eb",x"c2",x"87"),
  2595 => (x"74",x"78",x"c0",x"48"),
  2596 => (x"05",x"99",x"c8",x"49"),
  2597 => (x"f5",x"c3",x"87",x"ce"),
  2598 => (x"87",x"c7",x"e1",x"49"),
  2599 => (x"99",x"c2",x"49",x"70"),
  2600 => (x"87",x"ee",x"c0",x"02"),
  2601 => (x"bf",x"f6",x"c0",x"c3"),
  2602 => (x"87",x"c9",x"c0",x"02"),
  2603 => (x"c3",x"88",x"c1",x"48"),
  2604 => (x"d8",x"58",x"fa",x"c0"),
  2605 => (x"f2",x"c0",x"c3",x"87"),
  2606 => (x"91",x"cc",x"49",x"bf"),
  2607 => (x"c8",x"81",x"66",x"c4"),
  2608 => (x"bf",x"6e",x"7e",x"a1"),
  2609 => (x"87",x"c5",x"c0",x"02"),
  2610 => (x"73",x"49",x"ff",x"4b"),
  2611 => (x"48",x"a6",x"c8",x"0f"),
  2612 => (x"49",x"74",x"78",x"c1"),
  2613 => (x"c0",x"05",x"99",x"c4"),
  2614 => (x"f2",x"c3",x"87",x"ce"),
  2615 => (x"87",x"c3",x"e0",x"49"),
  2616 => (x"99",x"c2",x"49",x"70"),
  2617 => (x"87",x"fe",x"c0",x"02"),
  2618 => (x"c3",x"48",x"a6",x"c8"),
  2619 => (x"78",x"bf",x"f2",x"c0"),
  2620 => (x"c1",x"49",x"66",x"c8"),
  2621 => (x"f6",x"c0",x"c3",x"89"),
  2622 => (x"b7",x"6e",x"7e",x"bf"),
  2623 => (x"ca",x"c0",x"06",x"a9"),
  2624 => (x"80",x"c1",x"48",x"87"),
  2625 => (x"58",x"fa",x"c0",x"c3"),
  2626 => (x"c8",x"87",x"d6",x"c0"),
  2627 => (x"91",x"cc",x"49",x"66"),
  2628 => (x"c8",x"81",x"66",x"c4"),
  2629 => (x"bf",x"6e",x"7e",x"a1"),
  2630 => (x"87",x"c5",x"c0",x"02"),
  2631 => (x"73",x"49",x"fe",x"4b"),
  2632 => (x"48",x"a6",x"c8",x"0f"),
  2633 => (x"fd",x"c3",x"78",x"c1"),
  2634 => (x"f6",x"de",x"ff",x"49"),
  2635 => (x"c2",x"49",x"70",x"87"),
  2636 => (x"ee",x"c0",x"02",x"99"),
  2637 => (x"f6",x"c0",x"c3",x"87"),
  2638 => (x"c9",x"c0",x"02",x"bf"),
  2639 => (x"f6",x"c0",x"c3",x"87"),
  2640 => (x"c0",x"78",x"c0",x"48"),
  2641 => (x"c0",x"c3",x"87",x"d8"),
  2642 => (x"cc",x"49",x"bf",x"f2"),
  2643 => (x"81",x"66",x"c4",x"91"),
  2644 => (x"6e",x"7e",x"a1",x"c8"),
  2645 => (x"c5",x"c0",x"02",x"bf"),
  2646 => (x"49",x"fd",x"4b",x"87"),
  2647 => (x"a6",x"c8",x"0f",x"73"),
  2648 => (x"c3",x"78",x"c1",x"48"),
  2649 => (x"dd",x"ff",x"49",x"fa"),
  2650 => (x"49",x"70",x"87",x"f9"),
  2651 => (x"c1",x"02",x"99",x"c2"),
  2652 => (x"a6",x"c8",x"87",x"c0"),
  2653 => (x"f2",x"c0",x"c3",x"48"),
  2654 => (x"66",x"c8",x"78",x"bf"),
  2655 => (x"c4",x"88",x"c1",x"48"),
  2656 => (x"c0",x"c3",x"58",x"a6"),
  2657 => (x"6e",x"48",x"bf",x"f6"),
  2658 => (x"c0",x"03",x"a8",x"b7"),
  2659 => (x"c0",x"c3",x"87",x"c9"),
  2660 => (x"78",x"6e",x"48",x"f6"),
  2661 => (x"c8",x"87",x"d6",x"c0"),
  2662 => (x"91",x"cc",x"49",x"66"),
  2663 => (x"c8",x"81",x"66",x"c4"),
  2664 => (x"bf",x"6e",x"7e",x"a1"),
  2665 => (x"87",x"c5",x"c0",x"02"),
  2666 => (x"73",x"49",x"fc",x"4b"),
  2667 => (x"48",x"a6",x"c8",x"0f"),
  2668 => (x"c0",x"c3",x"78",x"c1"),
  2669 => (x"c0",x"4b",x"bf",x"f6"),
  2670 => (x"c0",x"06",x"ab",x"b7"),
  2671 => (x"8b",x"c1",x"87",x"c9"),
  2672 => (x"01",x"ab",x"b7",x"c0"),
  2673 => (x"74",x"87",x"f7",x"ff"),
  2674 => (x"99",x"f0",x"c3",x"49"),
  2675 => (x"87",x"cf",x"c0",x"05"),
  2676 => (x"ff",x"49",x"da",x"c1"),
  2677 => (x"70",x"87",x"cc",x"dc"),
  2678 => (x"02",x"99",x"c2",x"49"),
  2679 => (x"c3",x"87",x"e8",x"c2"),
  2680 => (x"7e",x"bf",x"ee",x"c0"),
  2681 => (x"bf",x"f6",x"c0",x"c3"),
  2682 => (x"ab",x"b7",x"c0",x"4b"),
  2683 => (x"87",x"d0",x"c0",x"06"),
  2684 => (x"80",x"cc",x"48",x"6e"),
  2685 => (x"c1",x"58",x"a6",x"c4"),
  2686 => (x"ab",x"b7",x"c0",x"8b"),
  2687 => (x"87",x"f0",x"ff",x"01"),
  2688 => (x"4a",x"bf",x"97",x"6e"),
  2689 => (x"c0",x"02",x"8a",x"c1"),
  2690 => (x"02",x"8a",x"87",x"f7"),
  2691 => (x"8a",x"87",x"d6",x"c0"),
  2692 => (x"87",x"ca",x"c1",x"02"),
  2693 => (x"ee",x"c1",x"05",x"8a"),
  2694 => (x"c8",x"4a",x"6e",x"87"),
  2695 => (x"f4",x"49",x"6a",x"82"),
  2696 => (x"e2",x"c1",x"87",x"eb"),
  2697 => (x"c8",x"4b",x"6e",x"87"),
  2698 => (x"c2",x"1e",x"6b",x"83"),
  2699 => (x"fd",x"1e",x"c0",x"dd"),
  2700 => (x"c8",x"87",x"c9",x"d9"),
  2701 => (x"c3",x"4b",x"6b",x"86"),
  2702 => (x"49",x"bf",x"f6",x"c0"),
  2703 => (x"c6",x"c1",x"0f",x"73"),
  2704 => (x"c8",x"49",x"6e",x"87"),
  2705 => (x"69",x"48",x"c1",x"81"),
  2706 => (x"c3",x"49",x"70",x"30"),
  2707 => (x"48",x"bf",x"ea",x"c0"),
  2708 => (x"c0",x"c3",x"b8",x"71"),
  2709 => (x"a6",x"c8",x"58",x"ee"),
  2710 => (x"c0",x"78",x"c1",x"48"),
  2711 => (x"49",x"6e",x"87",x"e9"),
  2712 => (x"48",x"6e",x"81",x"c8"),
  2713 => (x"a6",x"c8",x"80",x"cb"),
  2714 => (x"97",x"66",x"c4",x"58"),
  2715 => (x"a2",x"c1",x"4a",x"bf"),
  2716 => (x"49",x"69",x"97",x"4b"),
  2717 => (x"c0",x"04",x"ab",x"b7"),
  2718 => (x"4b",x"c0",x"87",x"c2"),
  2719 => (x"97",x"0b",x"66",x"c4"),
  2720 => (x"a6",x"c8",x"0b",x"7b"),
  2721 => (x"75",x"78",x"c1",x"48"),
  2722 => (x"e9",x"c0",x"02",x"9d"),
  2723 => (x"c0",x"02",x"6d",x"87"),
  2724 => (x"49",x"6d",x"87",x"e4"),
  2725 => (x"87",x"cb",x"d9",x"ff"),
  2726 => (x"99",x"c1",x"49",x"70"),
  2727 => (x"87",x"cb",x"c0",x"02"),
  2728 => (x"c3",x"4b",x"a5",x"c4"),
  2729 => (x"49",x"bf",x"f6",x"c0"),
  2730 => (x"c8",x"0f",x"4b",x"6b"),
  2731 => (x"c5",x"c0",x"02",x"85"),
  2732 => (x"ff",x"05",x"6d",x"87"),
  2733 => (x"66",x"c8",x"87",x"dc"),
  2734 => (x"87",x"c8",x"c0",x"02"),
  2735 => (x"bf",x"f6",x"c0",x"c3"),
  2736 => (x"87",x"fe",x"ee",x"49"),
  2737 => (x"cc",x"f1",x"8e",x"f4"),
  2738 => (x"11",x"12",x"58",x"87"),
  2739 => (x"1c",x"1b",x"1d",x"14"),
  2740 => (x"91",x"59",x"5a",x"23"),
  2741 => (x"eb",x"f2",x"f5",x"94"),
  2742 => (x"00",x"00",x"00",x"f4"),
  2743 => (x"00",x"00",x"00",x"00"),
  2744 => (x"00",x"00",x"00",x"00"),
  2745 => (x"14",x"12",x"58",x"00"),
  2746 => (x"1c",x"1b",x"1d",x"11"),
  2747 => (x"94",x"59",x"5a",x"23"),
  2748 => (x"eb",x"f2",x"f5",x"91"),
  2749 => (x"00",x"00",x"00",x"f4"),
  2750 => (x"00",x"00",x"2a",x"fc"),
  2751 => (x"50",x"50",x"55",x"53"),
  2752 => (x"20",x"54",x"52",x"4f"),
  2753 => (x"00",x"53",x"45",x"4e"),
  2754 => (x"00",x"00",x"1e",x"58"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

