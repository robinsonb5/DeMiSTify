library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e0c1c387",
    12 => x"86c0d04e",
    13 => x"49e0c1c3",
    14 => x"48ececc2",
    15 => x"0389d089",
    16 => x"404040c0",
    17 => x"d087f640",
    18 => x"50c00581",
    19 => x"f90589c1",
    20 => x"ececc287",
    21 => x"e8ecc24d",
    22 => x"02ad744c",
    23 => x"0f2487c4",
    24 => x"f3c187f7",
    25 => x"ecc287f5",
    26 => x"ecc24dec",
    27 => x"ad744cec",
    28 => x"c487c602",
    29 => x"f50f6c8c",
    30 => x"87fd0087",
    31 => x"5c5b5e0e",
    32 => x"86f00e5d",
    33 => x"a6c44cc0",
    34 => x"c078c048",
    35 => x"c04ba6e4",
    36 => x"484966e0",
    37 => x"e4c080c1",
    38 => x"481158a6",
    39 => x"7058a6c4",
    40 => x"f6c30298",
    41 => x"0266c487",
    42 => x"c487c6c3",
    43 => x"78c048a6",
    44 => x"f0c04a6e",
    45 => x"dac2028a",
    46 => x"8af3c087",
    47 => x"87dbc202",
    48 => x"dc028ac1",
    49 => x"028ac887",
    50 => x"c487c8c2",
    51 => x"87d1028a",
    52 => x"c1028ac3",
    53 => x"8ac287eb",
    54 => x"c387c602",
    55 => x"c9c2058a",
    56 => x"7383c487",
    57 => x"6989c449",
    58 => x"c1026e7e",
    59 => x"a6c887c8",
    60 => x"c478c048",
    61 => x"cc78c080",
    62 => x"4a6e4d66",
    63 => x"cf2ab7dc",
    64 => x"c4486e9a",
    65 => x"7258a630",
    66 => x"87c5029a",
    67 => x"c148a6c8",
    68 => x"06aac978",
    69 => x"f7c087c5",
    70 => x"c087c382",
    71 => x"66c882f0",
    72 => x"7287c702",
    73 => x"87f3c249",
    74 => x"85c184c1",
    75 => x"04adb7c8",
    76 => x"c187c7ff",
    77 => x"f0c087cf",
    78 => x"87dfc249",
    79 => x"c4c184c1",
    80 => x"7383c487",
    81 => x"6a8ac44a",
    82 => x"87dbc149",
    83 => x"4ca44970",
    84 => x"c487f2c0",
    85 => x"78c148a6",
    86 => x"c487eac0",
    87 => x"c44a7383",
    88 => x"c1496a8a",
    89 => x"84c187f5",
    90 => x"496e87db",
    91 => x"d487ecc1",
    92 => x"c0486e87",
    93 => x"c705a8e5",
    94 => x"48a6c487",
    95 => x"87c578c1",
    96 => x"d6c1496e",
    97 => x"66e0c087",
    98 => x"80c14849",
    99 => x"58a6e4c0",
   100 => x"a6c44811",
   101 => x"05987058",
   102 => x"7487cafc",
   103 => x"268ef048",
   104 => x"264c264d",
   105 => x"0e4f264b",
   106 => x"0e5c5b5e",
   107 => x"4cc04b71",
   108 => x"029a4a13",
   109 => x"497287cd",
   110 => x"c187e0c0",
   111 => x"9a4a1384",
   112 => x"7487f305",
   113 => x"264c2648",
   114 => x"1e4f264b",
   115 => x"73814873",
   116 => x"87c502a9",
   117 => x"f6055312",
   118 => x"1e4f2687",
   119 => x"4ac0ff1e",
   120 => x"c0c4486a",
   121 => x"58a6c498",
   122 => x"f3029870",
   123 => x"487a7187",
   124 => x"1e4f2626",
   125 => x"d4ff1e73",
   126 => x"7bffc34b",
   127 => x"ffc34a6b",
   128 => x"c8496b7b",
   129 => x"c3b17232",
   130 => x"4a6b7bff",
   131 => x"b27131c8",
   132 => x"6b7bffc3",
   133 => x"7232c849",
   134 => x"c44871b1",
   135 => x"264d2687",
   136 => x"264b264c",
   137 => x"5b5e0e4f",
   138 => x"710e5d5c",
   139 => x"4cd4ff4a",
   140 => x"ffc34872",
   141 => x"c27c7098",
   142 => x"05bfecec",
   143 => x"66d087c8",
   144 => x"d430c948",
   145 => x"66d058a6",
   146 => x"7129d849",
   147 => x"98ffc348",
   148 => x"66d07c70",
   149 => x"7129d049",
   150 => x"98ffc348",
   151 => x"66d07c70",
   152 => x"7129c849",
   153 => x"98ffc348",
   154 => x"66d07c70",
   155 => x"98ffc348",
   156 => x"49727c70",
   157 => x"487129d0",
   158 => x"7098ffc3",
   159 => x"c94b6c7c",
   160 => x"c34dfff0",
   161 => x"d005abff",
   162 => x"7cffc387",
   163 => x"8dc14b6c",
   164 => x"c387c602",
   165 => x"f002abff",
   166 => x"fd487387",
   167 => x"c01e87ff",
   168 => x"48d4ff49",
   169 => x"c178ffc3",
   170 => x"b7c8c381",
   171 => x"87f104a9",
   172 => x"731e4f26",
   173 => x"c487e71e",
   174 => x"c04bdff8",
   175 => x"f0ffc01e",
   176 => x"fd49f7c1",
   177 => x"86c487df",
   178 => x"c005a8c1",
   179 => x"d4ff87ea",
   180 => x"78ffc348",
   181 => x"c0c0c0c1",
   182 => x"c01ec0c0",
   183 => x"e9c1f0e1",
   184 => x"87c1fd49",
   185 => x"987086c4",
   186 => x"ff87ca05",
   187 => x"ffc348d4",
   188 => x"cb48c178",
   189 => x"87e6fe87",
   190 => x"fe058bc1",
   191 => x"48c087fd",
   192 => x"1e87defc",
   193 => x"d4ff1e73",
   194 => x"78ffc348",
   195 => x"fa49fecc",
   196 => x"4bd387d5",
   197 => x"ffc01ec0",
   198 => x"49c1c1f0",
   199 => x"c487c6fc",
   200 => x"05987086",
   201 => x"d4ff87ca",
   202 => x"78ffc348",
   203 => x"87cb48c1",
   204 => x"c187ebfd",
   205 => x"dbff058b",
   206 => x"fb48c087",
   207 => x"4d4387e3",
   208 => x"4d430044",
   209 => x"20383544",
   210 => x"200a6425",
   211 => x"4d430020",
   212 => x"5f383544",
   213 => x"64252032",
   214 => x"0020200a",
   215 => x"35444d43",
   216 => x"64252038",
   217 => x"0020200a",
   218 => x"43484453",
   219 => x"696e4920",
   220 => x"6c616974",
   221 => x"74617a69",
   222 => x"206e6f69",
   223 => x"6f727265",
   224 => x"000a2172",
   225 => x"5f646d63",
   226 => x"38444d43",
   227 => x"73657220",
   228 => x"736e6f70",
   229 => x"25203a65",
   230 => x"49000a64",
   231 => x"00525245",
   232 => x"00495053",
   233 => x"63204453",
   234 => x"20647261",
   235 => x"657a6973",
   236 => x"20736920",
   237 => x"000a6425",
   238 => x"74697257",
   239 => x"61662065",
   240 => x"64656c69",
   241 => x"5f63000a",
   242 => x"657a6973",
   243 => x"6c756d5f",
   244 => x"25203a74",
   245 => x"72202c64",
   246 => x"5f646165",
   247 => x"6c5f6c62",
   248 => x"203a6e65",
   249 => x"202c6425",
   250 => x"7a697363",
   251 => x"25203a65",
   252 => x"4d000a64",
   253 => x"20746c75",
   254 => x"000a6425",
   255 => x"62206425",
   256 => x"6b636f6c",
   257 => x"666f2073",
   258 => x"7a697320",
   259 => x"64252065",
   260 => x"6425000a",
   261 => x"6f6c6220",
   262 => x"20736b63",
   263 => x"3520666f",
   264 => x"62203231",
   265 => x"73657479",
   266 => x"5e0e000a",
   267 => x"0e5d5c5b",
   268 => x"f94dd4ff",
   269 => x"eac687e8",
   270 => x"f0e1c01e",
   271 => x"f749c8c1",
   272 => x"4b7087e3",
   273 => x"1ec4ce1e",
   274 => x"cc87f1f0",
   275 => x"02abc186",
   276 => x"eefa87c8",
   277 => x"c248c087",
   278 => x"d6f687ca",
   279 => x"cf497087",
   280 => x"c699ffff",
   281 => x"c802a9ea",
   282 => x"87d7fa87",
   283 => x"f3c148c0",
   284 => x"7dffc387",
   285 => x"f84cf1c0",
   286 => x"987087f8",
   287 => x"87cbc102",
   288 => x"ffc01ec0",
   289 => x"49fac1f0",
   290 => x"c487daf6",
   291 => x"9b4b7086",
   292 => x"87edc005",
   293 => x"1ec2cd1e",
   294 => x"c387e1ef",
   295 => x"4b6d7dff",
   296 => x"1ececd1e",
   297 => x"d087d5ef",
   298 => x"7dffc386",
   299 => x"737d7d7d",
   300 => x"99c0c149",
   301 => x"c187c502",
   302 => x"87e8c048",
   303 => x"e3c048c0",
   304 => x"cd1e7387",
   305 => x"f3ee1edc",
   306 => x"c286c887",
   307 => x"87cc05ac",
   308 => x"ee1ee8cd",
   309 => x"86c487e6",
   310 => x"87c848c0",
   311 => x"fe058cc1",
   312 => x"48c087d5",
   313 => x"0e87f6f4",
   314 => x"5d5c5b5e",
   315 => x"d0ff1e0e",
   316 => x"c0c0c84d",
   317 => x"ececc24b",
   318 => x"ce78c148",
   319 => x"e6f249e0",
   320 => x"6d4cc787",
   321 => x"c4987348",
   322 => x"987058a6",
   323 => x"6d87cc02",
   324 => x"c4987348",
   325 => x"987058a6",
   326 => x"c287f405",
   327 => x"87fef57d",
   328 => x"9873486d",
   329 => x"7058a6c4",
   330 => x"87cc0298",
   331 => x"9873486d",
   332 => x"7058a6c4",
   333 => x"87f40598",
   334 => x"1ec07dc3",
   335 => x"c1d0e5c0",
   336 => x"e0f349c0",
   337 => x"c186c487",
   338 => x"87c105a8",
   339 => x"05acc24c",
   340 => x"dbce87cb",
   341 => x"87cff149",
   342 => x"d8c148c0",
   343 => x"058cc187",
   344 => x"fb87e0fe",
   345 => x"ecc287c4",
   346 => x"987058f0",
   347 => x"c187cd05",
   348 => x"f0ffc01e",
   349 => x"f249d0c1",
   350 => x"86c487eb",
   351 => x"c348d4ff",
   352 => x"e7c578ff",
   353 => x"f4ecc287",
   354 => x"ce1e7058",
   355 => x"ebeb1ee4",
   356 => x"6d86c887",
   357 => x"c4987348",
   358 => x"987058a6",
   359 => x"6d87cc02",
   360 => x"c4987348",
   361 => x"987058a6",
   362 => x"c287f405",
   363 => x"48d4ff7d",
   364 => x"c178ffc3",
   365 => x"e4f12648",
   366 => x"5b5e0e87",
   367 => x"1e0e5d5c",
   368 => x"4bc0c0c8",
   369 => x"eec54cc0",
   370 => x"c44adfcd",
   371 => x"d4ff5ca6",
   372 => x"7cffc34c",
   373 => x"fec3486c",
   374 => x"c0c205a8",
   375 => x"05997187",
   376 => x"ff87e2c0",
   377 => x"7348bfd0",
   378 => x"58a6c498",
   379 => x"ce029870",
   380 => x"bfd0ff87",
   381 => x"c4987348",
   382 => x"987058a6",
   383 => x"ff87f205",
   384 => x"d1c448d0",
   385 => x"4866d478",
   386 => x"06a8b7c0",
   387 => x"c387e0c0",
   388 => x"4a6c7cff",
   389 => x"c7029971",
   390 => x"970a7187",
   391 => x"81c10a7a",
   392 => x"c14866d4",
   393 => x"58a6d888",
   394 => x"01a8b7c0",
   395 => x"c387e0ff",
   396 => x"717c7cff",
   397 => x"e1c00599",
   398 => x"bfd0ff87",
   399 => x"c4987348",
   400 => x"987058a6",
   401 => x"ff87ce02",
   402 => x"7348bfd0",
   403 => x"58a6c498",
   404 => x"f2059870",
   405 => x"48d0ff87",
   406 => x"4ac178d0",
   407 => x"058ac17e",
   408 => x"6e87eefd",
   409 => x"f4ee2648",
   410 => x"5b5e0e87",
   411 => x"711e0e5c",
   412 => x"c0c0c84a",
   413 => x"ff4cc04b",
   414 => x"ffc348d4",
   415 => x"bfd0ff78",
   416 => x"c4987348",
   417 => x"987058a6",
   418 => x"ff87ce02",
   419 => x"7348bfd0",
   420 => x"58a6c498",
   421 => x"f2059870",
   422 => x"48d0ff87",
   423 => x"ff78c3c4",
   424 => x"ffc348d4",
   425 => x"c01e7278",
   426 => x"d1c1f0ff",
   427 => x"87f5ed49",
   428 => x"987086c4",
   429 => x"87eec005",
   430 => x"d41ec0c8",
   431 => x"f8fb4966",
   432 => x"7086c487",
   433 => x"bfd0ff4c",
   434 => x"c4987348",
   435 => x"987058a6",
   436 => x"ff87ce02",
   437 => x"7348bfd0",
   438 => x"58a6c498",
   439 => x"f2059870",
   440 => x"48d0ff87",
   441 => x"487478c2",
   442 => x"87f3ec26",
   443 => x"5c5b5e0e",
   444 => x"c01e0e5d",
   445 => x"f0ffc01e",
   446 => x"ec49c9c1",
   447 => x"1ed287e7",
   448 => x"49faecc2",
   449 => x"c887f2fa",
   450 => x"c14dc086",
   451 => x"adb7d285",
   452 => x"c287f804",
   453 => x"bf97faec",
   454 => x"99c0c349",
   455 => x"05a9c0c1",
   456 => x"c287e7c0",
   457 => x"bf97c1ed",
   458 => x"c231d049",
   459 => x"bf97c2ed",
   460 => x"7232c84a",
   461 => x"c3edc2b1",
   462 => x"b14abf97",
   463 => x"ffcf4d71",
   464 => x"c19dffff",
   465 => x"c235ca85",
   466 => x"edc287de",
   467 => x"4bbf97c3",
   468 => x"9bc633c1",
   469 => x"97c4edc2",
   470 => x"b7c749bf",
   471 => x"c2b37129",
   472 => x"bf97ffec",
   473 => x"98cf4849",
   474 => x"c258a6c4",
   475 => x"bf97c0ed",
   476 => x"ca9cc34c",
   477 => x"c1edc234",
   478 => x"c249bf97",
   479 => x"c2b47131",
   480 => x"bf97c2ed",
   481 => x"99c0c349",
   482 => x"7129b7c6",
   483 => x"701e74b4",
   484 => x"cf1e731e",
   485 => x"e3e31ec6",
   486 => x"c183c287",
   487 => x"70307348",
   488 => x"f3cf1e4b",
   489 => x"87d4e31e",
   490 => x"66d848c1",
   491 => x"58a6dc30",
   492 => x"4d49a4c1",
   493 => x"1e709573",
   494 => x"fccf1e75",
   495 => x"87fce21e",
   496 => x"6e86e4c0",
   497 => x"b7c0c848",
   498 => x"87d206a8",
   499 => x"486e35c1",
   500 => x"c428b7c1",
   501 => x"c0c858a6",
   502 => x"ff01a8b7",
   503 => x"1e7587ee",
   504 => x"e21ed2d0",
   505 => x"86c887d6",
   506 => x"e8264875",
   507 => x"5e0e87ef",
   508 => x"710e5c5b",
   509 => x"d04cc04b",
   510 => x"b7c04866",
   511 => x"e3c006a8",
   512 => x"cc4a1387",
   513 => x"49bf9766",
   514 => x"c14866cc",
   515 => x"58a6d080",
   516 => x"02aab771",
   517 => x"48c187c4",
   518 => x"84c187cc",
   519 => x"acb766d0",
   520 => x"87ddff04",
   521 => x"87c248c0",
   522 => x"4c264d26",
   523 => x"4f264b26",
   524 => x"5c5b5e0e",
   525 => x"f5c20e5d",
   526 => x"78c048e0",
   527 => x"49ddefc0",
   528 => x"c287e4e5",
   529 => x"c01ed8ed",
   530 => x"87ddf849",
   531 => x"987086c4",
   532 => x"c087cc05",
   533 => x"e549c9ec",
   534 => x"48c087cd",
   535 => x"c087e7ca",
   536 => x"e549eaef",
   537 => x"4bc087c1",
   538 => x"48d8fac2",
   539 => x"1ec878c1",
   540 => x"1ec1f0c0",
   541 => x"49ceeec2",
   542 => x"c887f3fd",
   543 => x"05987086",
   544 => x"fac287c6",
   545 => x"78c048d8",
   546 => x"f0c01ec8",
   547 => x"eec21eca",
   548 => x"d9fd49ea",
   549 => x"7086c887",
   550 => x"87c60598",
   551 => x"48d8fac2",
   552 => x"fac278c0",
   553 => x"c01ebfd8",
   554 => x"ff1ed3f0",
   555 => x"c887cddf",
   556 => x"d8fac286",
   557 => x"f7c102bf",
   558 => x"d6f5c287",
   559 => x"1e49bf9f",
   560 => x"49d6f5c2",
   561 => x"a0c2f848",
   562 => x"d01e7189",
   563 => x"1ec0c81e",
   564 => x"1efbecc0",
   565 => x"87e4deff",
   566 => x"f4c286d4",
   567 => x"c24bbfde",
   568 => x"bf9fd6f5",
   569 => x"ead6c54a",
   570 => x"c8c005aa",
   571 => x"def4c287",
   572 => x"d4c04bbf",
   573 => x"d5e9ca87",
   574 => x"ccc002aa",
   575 => x"ddecc087",
   576 => x"87e3e249",
   577 => x"fdc748c0",
   578 => x"c01e7387",
   579 => x"ff1ef8ed",
   580 => x"c287e9dd",
   581 => x"731ed8ed",
   582 => x"87cdf549",
   583 => x"987086cc",
   584 => x"87c5c005",
   585 => x"ddc748c0",
   586 => x"d0eec087",
   587 => x"87f7e149",
   588 => x"1ee6f0c0",
   589 => x"87c4ddff",
   590 => x"f0c01ec8",
   591 => x"eec21efe",
   592 => x"e9fa49ea",
   593 => x"7086cc87",
   594 => x"c9c00598",
   595 => x"e0f5c287",
   596 => x"c078c148",
   597 => x"1ec887e4",
   598 => x"1ec7f1c0",
   599 => x"49ceeec2",
   600 => x"c887cbfa",
   601 => x"02987086",
   602 => x"c087cfc0",
   603 => x"ff1ef7ee",
   604 => x"c487c9dc",
   605 => x"c648c086",
   606 => x"f5c287cc",
   607 => x"49bf97d6",
   608 => x"05a9d5c1",
   609 => x"c287cdc0",
   610 => x"bf97d7f5",
   611 => x"a9eac249",
   612 => x"87c5c002",
   613 => x"edc548c0",
   614 => x"d8edc287",
   615 => x"c34cbf97",
   616 => x"c002ace9",
   617 => x"ebc387cc",
   618 => x"c5c002ac",
   619 => x"c548c087",
   620 => x"edc287d4",
   621 => x"49bf97e3",
   622 => x"ccc00599",
   623 => x"e4edc287",
   624 => x"c249bf97",
   625 => x"c5c002a9",
   626 => x"c448c087",
   627 => x"edc287f8",
   628 => x"48bf97e5",
   629 => x"58dcf5c2",
   630 => x"c14a4970",
   631 => x"e0f5c28a",
   632 => x"711e725a",
   633 => x"d0f1c01e",
   634 => x"cfdaff1e",
   635 => x"c286cc87",
   636 => x"bf97e6ed",
   637 => x"c2817349",
   638 => x"bf97e7ed",
   639 => x"35c84d4a",
   640 => x"f9c28571",
   641 => x"edc25df8",
   642 => x"48bf97e8",
   643 => x"58ccfac2",
   644 => x"bfe0f5c2",
   645 => x"87dcc202",
   646 => x"efc01ec8",
   647 => x"eec21ed4",
   648 => x"c9f749ea",
   649 => x"7086c887",
   650 => x"c5c00298",
   651 => x"c348c087",
   652 => x"f5c287d4",
   653 => x"484abfd8",
   654 => x"f5c230c4",
   655 => x"fac258e8",
   656 => x"edc25ac8",
   657 => x"49bf97fd",
   658 => x"edc231c8",
   659 => x"4bbf97fc",
   660 => x"edc249a1",
   661 => x"4bbf97fe",
   662 => x"a17333d0",
   663 => x"ffedc249",
   664 => x"d84bbf97",
   665 => x"49a17333",
   666 => x"59d0fac2",
   667 => x"bfc8fac2",
   668 => x"f4f9c291",
   669 => x"f9c281bf",
   670 => x"eec259fc",
   671 => x"4bbf97c5",
   672 => x"eec233c8",
   673 => x"4cbf97c4",
   674 => x"eec24ba3",
   675 => x"4cbf97c6",
   676 => x"a37434d0",
   677 => x"c7eec24b",
   678 => x"cf4cbf97",
   679 => x"7434d89c",
   680 => x"fac24ba3",
   681 => x"8bc25bc0",
   682 => x"fac29273",
   683 => x"a17248c0",
   684 => x"87cbc178",
   685 => x"97eaedc2",
   686 => x"31c849bf",
   687 => x"97e9edc2",
   688 => x"49a14abf",
   689 => x"59e8f5c2",
   690 => x"ffc731c5",
   691 => x"c229c981",
   692 => x"c259c8fa",
   693 => x"bf97efed",
   694 => x"c232c84a",
   695 => x"bf97eeed",
   696 => x"c24aa24b",
   697 => x"c25ad0fa",
   698 => x"92bfc8fa",
   699 => x"fac28275",
   700 => x"f9c25ac4",
   701 => x"78c048fc",
   702 => x"48f8f9c2",
   703 => x"c078a172",
   704 => x"87e3cd49",
   705 => x"dff448c1",
   706 => x"61655287",
   707 => x"666f2064",
   708 => x"52424d20",
   709 => x"69616620",
   710 => x"0a64656c",
   711 => x"206f4e00",
   712 => x"74726170",
   713 => x"6f697469",
   714 => x"6973206e",
   715 => x"74616e67",
   716 => x"20657275",
   717 => x"6e756f66",
   718 => x"4d000a64",
   719 => x"69735242",
   720 => x"203a657a",
   721 => x"202c6425",
   722 => x"74726170",
   723 => x"6f697469",
   724 => x"7a69736e",
   725 => x"25203a65",
   726 => x"6f202c64",
   727 => x"65736666",
   728 => x"666f2074",
   729 => x"67697320",
   730 => x"6425203a",
   731 => x"6973202c",
   732 => x"78302067",
   733 => x"000a7825",
   734 => x"64616552",
   735 => x"20676e69",
   736 => x"746f6f62",
   737 => x"63657320",
   738 => x"20726f74",
   739 => x"000a6425",
   740 => x"64616552",
   741 => x"6f6f6220",
   742 => x"65732074",
   743 => x"726f7463",
   744 => x"6f726620",
   745 => x"6966206d",
   746 => x"20747372",
   747 => x"74726170",
   748 => x"6f697469",
   749 => x"55000a6e",
   750 => x"7075736e",
   751 => x"74726f70",
   752 => x"70206465",
   753 => x"69747261",
   754 => x"6e6f6974",
   755 => x"70797420",
   756 => x"000d2165",
   757 => x"33544146",
   758 => x"20202032",
   759 => x"61655200",
   760 => x"676e6964",
   761 => x"52424d20",
   762 => x"424d000a",
   763 => x"75732052",
   764 => x"73656363",
   765 => x"6c756673",
   766 => x"7220796c",
   767 => x"0a646165",
   768 => x"54414600",
   769 => x"20203631",
   770 => x"41460020",
   771 => x"20323354",
   772 => x"50002020",
   773 => x"69747261",
   774 => x"6e6f6974",
   775 => x"6e756f63",
   776 => x"64252074",
   777 => x"7548000a",
   778 => x"6e69746e",
   779 => x"6f662067",
   780 => x"69662072",
   781 => x"7973656c",
   782 => x"6d657473",
   783 => x"4146000a",
   784 => x"20323354",
   785 => x"46002020",
   786 => x"36315441",
   787 => x"00202020",
   788 => x"73756c43",
   789 => x"20726574",
   790 => x"657a6973",
   791 => x"6425203a",
   792 => x"6c43202c",
   793 => x"65747375",
   794 => x"616d2072",
   795 => x"202c6b73",
   796 => x"000a6425",
   797 => x"6e65704f",
   798 => x"66206465",
   799 => x"2c656c69",
   800 => x"616f6c20",
   801 => x"676e6964",
   802 => x"0a2e2e2e",
   803 => x"6e614300",
   804 => x"6f207427",
   805 => x"206e6570",
   806 => x"000a7325",
   807 => x"5c5b5e0e",
   808 => x"4a710e5d",
   809 => x"bfe0f5c2",
   810 => x"7287cc02",
   811 => x"2bb7c74b",
   812 => x"ffc14d72",
   813 => x"7287ca9d",
   814 => x"2bb7c84b",
   815 => x"ffc34d72",
   816 => x"d8edc29d",
   817 => x"f4f9c21e",
   818 => x"817349bf",
   819 => x"87d9e671",
   820 => x"987086c4",
   821 => x"c087c505",
   822 => x"87e6c048",
   823 => x"bfe0f5c2",
   824 => x"7587d202",
   825 => x"c291c449",
   826 => x"6981d8ed",
   827 => x"ffffcf4c",
   828 => x"cb9cffff",
   829 => x"c2497587",
   830 => x"d8edc291",
   831 => x"4c699f81",
   832 => x"e3ec4874",
   833 => x"5b5e0e87",
   834 => x"f40e5d5c",
   835 => x"c04c7186",
   836 => x"d0fac24b",
   837 => x"a6c47ebf",
   838 => x"d4fac248",
   839 => x"a6c878bf",
   840 => x"c278c048",
   841 => x"48bfe4f5",
   842 => x"c206a8c0",
   843 => x"66c887e3",
   844 => x"0599cf49",
   845 => x"edc287d8",
   846 => x"66c81ed8",
   847 => x"80c14849",
   848 => x"e458a6cc",
   849 => x"86c487e3",
   850 => x"4bd8edc2",
   851 => x"e0c087c3",
   852 => x"4a6b9783",
   853 => x"e7c1029a",
   854 => x"aae5c387",
   855 => x"87e0c102",
   856 => x"9749a3cb",
   857 => x"99d84969",
   858 => x"87d4c105",
   859 => x"d0ff4973",
   860 => x"1ecb87f5",
   861 => x"1e66e0c0",
   862 => x"f1e94973",
   863 => x"7086c887",
   864 => x"fbc00598",
   865 => x"4aa3dc87",
   866 => x"6a49a4c4",
   867 => x"49a3da79",
   868 => x"9f4da4c8",
   869 => x"c27d4869",
   870 => x"02bfe0f5",
   871 => x"a3d487d3",
   872 => x"49699f49",
   873 => x"99ffffc0",
   874 => x"30d04871",
   875 => x"c258a6c4",
   876 => x"6e7ec087",
   877 => x"70806d48",
   878 => x"c17cc07d",
   879 => x"87c5c148",
   880 => x"c14866c8",
   881 => x"58a6cc80",
   882 => x"bfe4f5c2",
   883 => x"ddfd04a8",
   884 => x"e0f5c287",
   885 => x"eac002bf",
   886 => x"fa496e87",
   887 => x"a6c487fe",
   888 => x"cf497058",
   889 => x"f8ffffff",
   890 => x"d602a999",
   891 => x"c2497087",
   892 => x"d8f5c289",
   893 => x"f9c291bf",
   894 => x"7148bff8",
   895 => x"58a6c880",
   896 => x"c087dbfc",
   897 => x"e88ef448",
   898 => x"731e87de",
   899 => x"6a4a711e",
   900 => x"7181c149",
   901 => x"dcf5c27a",
   902 => x"cb0599bf",
   903 => x"4ba2c887",
   904 => x"f7f9496b",
   905 => x"7b497087",
   906 => x"ffe748c1",
   907 => x"1e731e87",
   908 => x"f9c24b71",
   909 => x"c849bff8",
   910 => x"4a6a4aa3",
   911 => x"f5c28ac2",
   912 => x"7292bfd8",
   913 => x"f5c249a1",
   914 => x"6b4abfdc",
   915 => x"49a1729a",
   916 => x"711e66c8",
   917 => x"c487d2e0",
   918 => x"05987086",
   919 => x"48c087c4",
   920 => x"48c187c2",
   921 => x"0e87c5e7",
   922 => x"0e5c5b5e",
   923 => x"4bc04a71",
   924 => x"c0029a72",
   925 => x"a2da87e0",
   926 => x"4b699f49",
   927 => x"bfe0f5c2",
   928 => x"d487cf02",
   929 => x"699f49a2",
   930 => x"ffc04c49",
   931 => x"34d09cff",
   932 => x"4cc087c2",
   933 => x"9b73b374",
   934 => x"4a87df02",
   935 => x"f5c28ac2",
   936 => x"9249bfd8",
   937 => x"bff8f9c2",
   938 => x"c2807248",
   939 => x"7158d8fa",
   940 => x"c230c448",
   941 => x"c058e8f5",
   942 => x"f9c287e9",
   943 => x"c24bbffc",
   944 => x"c248d4fa",
   945 => x"78bfc0fa",
   946 => x"bfe0f5c2",
   947 => x"c287c902",
   948 => x"49bfd8f5",
   949 => x"87c731c4",
   950 => x"bfc4fac2",
   951 => x"c231c449",
   952 => x"c259e8f5",
   953 => x"e55bd4fa",
   954 => x"5e0e87c0",
   955 => x"0e5d5c5b",
   956 => x"4a7186f4",
   957 => x"87de029a",
   958 => x"48d4edc2",
   959 => x"edc278c0",
   960 => x"fac248cc",
   961 => x"c278bfd4",
   962 => x"c248d0ed",
   963 => x"78bfd0fa",
   964 => x"48c2c3c1",
   965 => x"f5c278c0",
   966 => x"c249bfe4",
   967 => x"4abfd4ed",
   968 => x"c403aa71",
   969 => x"497287cc",
   970 => x"c00599cf",
   971 => x"edc287e1",
   972 => x"edc21ed8",
   973 => x"c249bfcc",
   974 => x"c148cced",
   975 => x"ff7178a1",
   976 => x"c487e6dc",
   977 => x"fec2c186",
   978 => x"d8edc248",
   979 => x"c187cc78",
   980 => x"48bffec2",
   981 => x"c180e0c0",
   982 => x"c258c2c3",
   983 => x"48bfd4ed",
   984 => x"edc280c1",
   985 => x"be2758d8",
   986 => x"bf000010",
   987 => x"9c4cbf97",
   988 => x"87eec202",
   989 => x"02ace5c3",
   990 => x"c187e7c2",
   991 => x"4bbffec2",
   992 => x"1149a3cb",
   993 => x"05adcf4d",
   994 => x"7487d6c1",
   995 => x"c199df49",
   996 => x"c291cd89",
   997 => x"c181e8f5",
   998 => x"51124aa3",
   999 => x"124aa3c3",
  1000 => x"4aa3c551",
  1001 => x"a3c75112",
  1002 => x"c951124a",
  1003 => x"51124aa3",
  1004 => x"124aa3ce",
  1005 => x"4aa3d051",
  1006 => x"a3d25112",
  1007 => x"d451124a",
  1008 => x"51124aa3",
  1009 => x"124aa3d6",
  1010 => x"4aa3d851",
  1011 => x"a3dc5112",
  1012 => x"de51124a",
  1013 => x"51124aa3",
  1014 => x"48c2c3c1",
  1015 => x"c1c178c1",
  1016 => x"c8497587",
  1017 => x"f3c00599",
  1018 => x"d0497587",
  1019 => x"87d00599",
  1020 => x"c00266dc",
  1021 => x"497387ca",
  1022 => x"700f66dc",
  1023 => x"87dc0298",
  1024 => x"bfc2c3c1",
  1025 => x"87c6c005",
  1026 => x"48e8f5c2",
  1027 => x"c3c150c0",
  1028 => x"78c048c2",
  1029 => x"bffec2c1",
  1030 => x"87dcc248",
  1031 => x"48c2c3c1",
  1032 => x"f5c278c0",
  1033 => x"c249bfe4",
  1034 => x"4abfd4ed",
  1035 => x"fb04aa71",
  1036 => x"fac287f4",
  1037 => x"c005bfd4",
  1038 => x"f5c287c8",
  1039 => x"c102bfe0",
  1040 => x"edc287f4",
  1041 => x"f149bfd0",
  1042 => x"edc287d2",
  1043 => x"7e7058d4",
  1044 => x"bfe0f5c2",
  1045 => x"87ddc002",
  1046 => x"ffcf496e",
  1047 => x"99f8ffff",
  1048 => x"c8c002a9",
  1049 => x"48a6c487",
  1050 => x"e6c078c0",
  1051 => x"48a6c487",
  1052 => x"dec078c1",
  1053 => x"cf496e87",
  1054 => x"a999f8ff",
  1055 => x"87c8c002",
  1056 => x"c048a6c8",
  1057 => x"87c5c078",
  1058 => x"c148a6c8",
  1059 => x"48a6c478",
  1060 => x"c47866c8",
  1061 => x"ddc00566",
  1062 => x"c2496e87",
  1063 => x"d8f5c289",
  1064 => x"f9c291bf",
  1065 => x"7148bff8",
  1066 => x"d0edc280",
  1067 => x"d4edc258",
  1068 => x"f978c048",
  1069 => x"48c087e0",
  1070 => x"ddff8ef4",
  1071 => x"000087ea",
  1072 => x"00000000",
  1073 => x"ff1e0000",
  1074 => x"ffc348d4",
  1075 => x"99496878",
  1076 => x"c087c602",
  1077 => x"ee05a9fb",
  1078 => x"26487187",
  1079 => x"5b5e0e4f",
  1080 => x"4a710e5c",
  1081 => x"d4ff4bc0",
  1082 => x"78ffc348",
  1083 => x"02994968",
  1084 => x"c087c1c1",
  1085 => x"c002a9ec",
  1086 => x"fbc087fa",
  1087 => x"f3c002a9",
  1088 => x"b766cc87",
  1089 => x"87cc03ab",
  1090 => x"c70266d0",
  1091 => x"97097287",
  1092 => x"82c10979",
  1093 => x"c2029971",
  1094 => x"ff83c187",
  1095 => x"ffc348d4",
  1096 => x"99496878",
  1097 => x"c087cd02",
  1098 => x"c702a9ec",
  1099 => x"a9fbc087",
  1100 => x"87cdff05",
  1101 => x"c30266d0",
  1102 => x"7a97c087",
  1103 => x"05a9fbc0",
  1104 => x"4c7387c7",
  1105 => x"c28c0cc0",
  1106 => x"744c7387",
  1107 => x"2687c248",
  1108 => x"264c264d",
  1109 => x"1e4f264b",
  1110 => x"c348d4ff",
  1111 => x"496878ff",
  1112 => x"a9b7f0c0",
  1113 => x"c087ca04",
  1114 => x"01a9b7f9",
  1115 => x"f0c087c3",
  1116 => x"b7c1c189",
  1117 => x"87ca04a9",
  1118 => x"a9b7c6c1",
  1119 => x"c087c301",
  1120 => x"487189f7",
  1121 => x"5e0e4f26",
  1122 => x"0e5d5c5b",
  1123 => x"4c7186f4",
  1124 => x"c04bd4ff",
  1125 => x"ffc37e4d",
  1126 => x"bfd0ff7b",
  1127 => x"c0c0c848",
  1128 => x"58a6c898",
  1129 => x"d0029870",
  1130 => x"bfd0ff87",
  1131 => x"c0c0c848",
  1132 => x"58a6c898",
  1133 => x"f0059870",
  1134 => x"48d0ff87",
  1135 => x"d478e1c0",
  1136 => x"87c2fc7b",
  1137 => x"02994970",
  1138 => x"c387c7c1",
  1139 => x"a6c87bff",
  1140 => x"c8786b48",
  1141 => x"fbc04866",
  1142 => x"87c802a8",
  1143 => x"bff0fac2",
  1144 => x"87eec002",
  1145 => x"99714dc1",
  1146 => x"87e6c002",
  1147 => x"02a9fbc0",
  1148 => x"d1fb87c3",
  1149 => x"7bffc387",
  1150 => x"c6c1496b",
  1151 => x"87cc05a9",
  1152 => x"7b7bffc3",
  1153 => x"6b48a6c8",
  1154 => x"4d49c078",
  1155 => x"ff059971",
  1156 => x"9d7587da",
  1157 => x"87dec105",
  1158 => x"6b7bffc3",
  1159 => x"7bffc34a",
  1160 => x"6b48a6c4",
  1161 => x"c1486e78",
  1162 => x"58a6c480",
  1163 => x"9749a4c8",
  1164 => x"66c84969",
  1165 => x"87da05a9",
  1166 => x"9749a4c9",
  1167 => x"05aa4969",
  1168 => x"a4ca87d0",
  1169 => x"49699749",
  1170 => x"05a966c4",
  1171 => x"4dc187c4",
  1172 => x"66c887d6",
  1173 => x"a8ecc048",
  1174 => x"c887c902",
  1175 => x"fbc04866",
  1176 => x"87c405a8",
  1177 => x"4dc17ec0",
  1178 => x"c87bffc3",
  1179 => x"786b48a6",
  1180 => x"fe029d75",
  1181 => x"d0ff87e2",
  1182 => x"c0c848bf",
  1183 => x"a6c898c0",
  1184 => x"02987058",
  1185 => x"d0ff87d0",
  1186 => x"c0c848bf",
  1187 => x"a6c898c0",
  1188 => x"05987058",
  1189 => x"d0ff87f0",
  1190 => x"78e0c048",
  1191 => x"8ef4486e",
  1192 => x"0e87ecfa",
  1193 => x"5d5c5b5e",
  1194 => x"c486f40e",
  1195 => x"d0ff59a6",
  1196 => x"c0c0c84c",
  1197 => x"c21e6e4b",
  1198 => x"e949f4fa",
  1199 => x"86c487c7",
  1200 => x"c6029870",
  1201 => x"fac287cb",
  1202 => x"6e4dbff8",
  1203 => x"87f6fa49",
  1204 => x"7058a6c8",
  1205 => x"4966c41e",
  1206 => x"1e7181c8",
  1207 => x"1ed8d1c1",
  1208 => x"87d8f6fe",
  1209 => x"486c86cc",
  1210 => x"a6cc9873",
  1211 => x"02987058",
  1212 => x"486c87cc",
  1213 => x"a6c49873",
  1214 => x"05987058",
  1215 => x"7cc587f4",
  1216 => x"c148d4ff",
  1217 => x"fac278d5",
  1218 => x"c149bff0",
  1219 => x"4a66c481",
  1220 => x"32c68ac1",
  1221 => x"b0714872",
  1222 => x"7808d4ff",
  1223 => x"9873486c",
  1224 => x"7058a6c4",
  1225 => x"87cc0298",
  1226 => x"9873486c",
  1227 => x"7058a6c4",
  1228 => x"87f40598",
  1229 => x"d4ff7cc4",
  1230 => x"78ffc348",
  1231 => x"9873486c",
  1232 => x"7058a6c4",
  1233 => x"87cc0298",
  1234 => x"9873486c",
  1235 => x"7058a6c4",
  1236 => x"87f40598",
  1237 => x"d4ff7cc5",
  1238 => x"78d3c148",
  1239 => x"486c78c1",
  1240 => x"a6c49873",
  1241 => x"02987058",
  1242 => x"486c87cc",
  1243 => x"a6c49873",
  1244 => x"05987058",
  1245 => x"7cc487f4",
  1246 => x"c2029d75",
  1247 => x"edc287d1",
  1248 => x"c21e7ed8",
  1249 => x"ea49f4fa",
  1250 => x"86c487e3",
  1251 => x"c5059870",
  1252 => x"c248c087",
  1253 => x"c0c887fd",
  1254 => x"c404adb7",
  1255 => x"c48d4a87",
  1256 => x"c04a7587",
  1257 => x"73486c4d",
  1258 => x"58a6c898",
  1259 => x"cc029870",
  1260 => x"73486c87",
  1261 => x"58a6c898",
  1262 => x"f4059870",
  1263 => x"ff7ccd87",
  1264 => x"d4c148d4",
  1265 => x"c1497278",
  1266 => x"0299718a",
  1267 => x"976e87d9",
  1268 => x"d4ff48bf",
  1269 => x"486e7808",
  1270 => x"a6c480c1",
  1271 => x"c1497258",
  1272 => x"0599718a",
  1273 => x"6c87e7ff",
  1274 => x"c4987348",
  1275 => x"987058a6",
  1276 => x"6c87cd02",
  1277 => x"c4987348",
  1278 => x"987058a6",
  1279 => x"87f3ff05",
  1280 => x"fac27cc4",
  1281 => x"c1e849f4",
  1282 => x"059d7587",
  1283 => x"6c87effd",
  1284 => x"c4987348",
  1285 => x"987058a6",
  1286 => x"6c87cd02",
  1287 => x"c4987348",
  1288 => x"987058a6",
  1289 => x"87f3ff05",
  1290 => x"d4ff7cc5",
  1291 => x"78d3c148",
  1292 => x"486c78c0",
  1293 => x"a6c49873",
  1294 => x"02987058",
  1295 => x"486c87cd",
  1296 => x"a6c49873",
  1297 => x"05987058",
  1298 => x"c487f3ff",
  1299 => x"c248c17c",
  1300 => x"f448c087",
  1301 => x"87f7f38e",
  1302 => x"6e65704f",
  1303 => x"66206465",
  1304 => x"2c656c69",
  1305 => x"616f6c20",
  1306 => x"676e6964",
  1307 => x"2c732520",
  1308 => x"64692820",
  1309 => x"64252078",
  1310 => x"2e2e2e29",
  1311 => x"6f4c000a",
  1312 => x"6e696461",
  1313 => x"2e2e2e67",
  1314 => x"6c694600",
  1315 => x"73252065",
  1316 => x"2080000a",
  1317 => x"6b636142",
  1318 => x"616f4c00",
  1319 => x"2e2a2064",
  1320 => x"203a0020",
  1321 => x"42208000",
  1322 => x"006b6361",
  1323 => x"78452080",
  1324 => x"49007469",
  1325 => x"6974696e",
  1326 => x"7a696c61",
  1327 => x"20676e69",
  1328 => x"63204453",
  1329 => x"0a647261",
  1330 => x"76614800",
  1331 => x"44532065",
  1332 => x"4f42000a",
  1333 => x"2020544f",
  1334 => x"4f522020",
  1335 => x"5e0e004d",
  1336 => x"0e5d5c5b",
  1337 => x"c04b711e",
  1338 => x"abb74d4c",
  1339 => x"87e9c004",
  1340 => x"1ec6c6c1",
  1341 => x"c4029d75",
  1342 => x"c24ac087",
  1343 => x"724ac187",
  1344 => x"87e6e749",
  1345 => x"58a686c4",
  1346 => x"056e84c1",
  1347 => x"4c7387c2",
  1348 => x"b77385c1",
  1349 => x"d7ff06ac",
  1350 => x"26486e87",
  1351 => x"0e87f0f0",
  1352 => x"5d5c5b5e",
  1353 => x"4c711e0e",
  1354 => x"c4fbc249",
  1355 => x"edfe81bf",
  1356 => x"1e4d7087",
  1357 => x"1ec9d2c1",
  1358 => x"87c0edfe",
  1359 => x"9d7586c8",
  1360 => x"87fcc002",
  1361 => x"4be8f5c2",
  1362 => x"49cb4a75",
  1363 => x"87fbf1fe",
  1364 => x"91de4974",
  1365 => x"48d8fbc2",
  1366 => x"a6c48071",
  1367 => x"fed1c158",
  1368 => x"c8496e48",
  1369 => x"41204aa1",
  1370 => x"f905aa71",
  1371 => x"10511087",
  1372 => x"74511051",
  1373 => x"e9c4c149",
  1374 => x"e8f5c287",
  1375 => x"87e3f449",
  1376 => x"49c4f7c1",
  1377 => x"87e5c7c1",
  1378 => x"87c1c8c1",
  1379 => x"87ffee26",
  1380 => x"711e731e",
  1381 => x"fbc2494b",
  1382 => x"fd81bfc4",
  1383 => x"4a7087c0",
  1384 => x"87c4029a",
  1385 => x"87ffe249",
  1386 => x"48c4fbc2",
  1387 => x"497378c0",
  1388 => x"ee87e9c1",
  1389 => x"731e87dd",
  1390 => x"c44b711e",
  1391 => x"c1024aa3",
  1392 => x"8ac187c8",
  1393 => x"8a87dc02",
  1394 => x"87f1c002",
  1395 => x"c4c1058a",
  1396 => x"c4fbc287",
  1397 => x"fcc002bf",
  1398 => x"88c14887",
  1399 => x"58c8fbc2",
  1400 => x"c287f2c0",
  1401 => x"49bfc4fb",
  1402 => x"fbc289d0",
  1403 => x"b7c059c8",
  1404 => x"e0c003a9",
  1405 => x"c4fbc287",
  1406 => x"d878c048",
  1407 => x"c4fbc287",
  1408 => x"80c148bf",
  1409 => x"58c8fbc2",
  1410 => x"fbc287cb",
  1411 => x"d048bfc4",
  1412 => x"c8fbc280",
  1413 => x"c3497358",
  1414 => x"87f7ec87",
  1415 => x"5c5b5e0e",
  1416 => x"86f00e5d",
  1417 => x"c259a6d0",
  1418 => x"c04dd8ed",
  1419 => x"48a6c44c",
  1420 => x"fbc278c0",
  1421 => x"c048bfc4",
  1422 => x"c106a8b7",
  1423 => x"edc287c1",
  1424 => x"029848d8",
  1425 => x"c187f8c0",
  1426 => x"c81ec6c6",
  1427 => x"87c70266",
  1428 => x"c048a6c4",
  1429 => x"c487c578",
  1430 => x"78c148a6",
  1431 => x"e24966c4",
  1432 => x"86c487c8",
  1433 => x"84c14d70",
  1434 => x"c14866c4",
  1435 => x"58a6c880",
  1436 => x"bfc4fbc2",
  1437 => x"c603acb7",
  1438 => x"059d7587",
  1439 => x"c087c8ff",
  1440 => x"029d754c",
  1441 => x"c187e3c3",
  1442 => x"c81ec6c6",
  1443 => x"87c70266",
  1444 => x"c048a6cc",
  1445 => x"cc87c578",
  1446 => x"78c148a6",
  1447 => x"e14966cc",
  1448 => x"86c487c8",
  1449 => x"026e58a6",
  1450 => x"4987ebc2",
  1451 => x"699781cb",
  1452 => x"0299d049",
  1453 => x"c187d9c1",
  1454 => x"744bd0d6",
  1455 => x"c191cc49",
  1456 => x"c881c4f7",
  1457 => x"7a734aa1",
  1458 => x"ffc381c1",
  1459 => x"de497451",
  1460 => x"d8fbc291",
  1461 => x"c285714d",
  1462 => x"c17d97c1",
  1463 => x"e0c049a5",
  1464 => x"e8f5c251",
  1465 => x"d202bf97",
  1466 => x"c284c187",
  1467 => x"f5c24ba5",
  1468 => x"49db4ae8",
  1469 => x"87d3ebfe",
  1470 => x"cd87dbc1",
  1471 => x"51c049a5",
  1472 => x"a5c284c1",
  1473 => x"cb4a6e4b",
  1474 => x"feeafe49",
  1475 => x"87c6c187",
  1476 => x"91cc4974",
  1477 => x"81c4f7c1",
  1478 => x"d4c181c8",
  1479 => x"f5c279df",
  1480 => x"02bf97e8",
  1481 => x"497487d8",
  1482 => x"84c191de",
  1483 => x"4bd8fbc2",
  1484 => x"f5c28371",
  1485 => x"49dd4ae8",
  1486 => x"87cfeafe",
  1487 => x"4b7487d8",
  1488 => x"fbc293de",
  1489 => x"a3cb83d8",
  1490 => x"c151c049",
  1491 => x"4a6e7384",
  1492 => x"e9fe49cb",
  1493 => x"66c487f5",
  1494 => x"c880c148",
  1495 => x"b7c758a6",
  1496 => x"c5c003ac",
  1497 => x"fc056e87",
  1498 => x"b7c787dd",
  1499 => x"d3c003ac",
  1500 => x"de497487",
  1501 => x"d8fbc291",
  1502 => x"c151c081",
  1503 => x"acb7c784",
  1504 => x"87edff04",
  1505 => x"48d9f8c1",
  1506 => x"f8c150c0",
  1507 => x"50c248d8",
  1508 => x"48e0f8c1",
  1509 => x"78c2dfc1",
  1510 => x"48dcf8c1",
  1511 => x"78d2d2c1",
  1512 => x"48ecf8c1",
  1513 => x"78f6d6c1",
  1514 => x"c04966cc",
  1515 => x"f087f3fb",
  1516 => x"87dbe68e",
  1517 => x"c24a711e",
  1518 => x"725af4fa",
  1519 => x"87dcf949",
  1520 => x"711e4f26",
  1521 => x"91cc494a",
  1522 => x"81c4f7c1",
  1523 => x"481181c1",
  1524 => x"58f0fac2",
  1525 => x"49a2f0c0",
  1526 => x"87ffe7fe",
  1527 => x"ddd549c0",
  1528 => x"0e4f2687",
  1529 => x"5d5c5b5e",
  1530 => x"7186f00e",
  1531 => x"91cc494c",
  1532 => x"81c4f7c1",
  1533 => x"c47ea1c3",
  1534 => x"fac248a6",
  1535 => x"6e78bfe8",
  1536 => x"c44abf97",
  1537 => x"2b724b66",
  1538 => x"124aa1c1",
  1539 => x"58a6cc48",
  1540 => x"83c19b70",
  1541 => x"699781c2",
  1542 => x"04abb749",
  1543 => x"4bc087c2",
  1544 => x"4abf976e",
  1545 => x"724966c8",
  1546 => x"c4b9ff31",
  1547 => x"4d739966",
  1548 => x"b5713572",
  1549 => x"5decfac2",
  1550 => x"c348d4ff",
  1551 => x"d0ff78ff",
  1552 => x"c0c848bf",
  1553 => x"a6d098c0",
  1554 => x"02987058",
  1555 => x"d0ff87d0",
  1556 => x"c0c848bf",
  1557 => x"a6c498c0",
  1558 => x"05987058",
  1559 => x"d0ff87f0",
  1560 => x"78e1c048",
  1561 => x"de48d4ff",
  1562 => x"7d0d7078",
  1563 => x"c848750d",
  1564 => x"d4ff28b7",
  1565 => x"48757808",
  1566 => x"ff28b7d0",
  1567 => x"757808d4",
  1568 => x"28b7d848",
  1569 => x"7808d4ff",
  1570 => x"48bfd0ff",
  1571 => x"98c0c0c8",
  1572 => x"7058a6c4",
  1573 => x"87d00298",
  1574 => x"48bfd0ff",
  1575 => x"98c0c0c8",
  1576 => x"7058a6c4",
  1577 => x"87f00598",
  1578 => x"c048d0ff",
  1579 => x"1ec778e0",
  1580 => x"f7c11ec0",
  1581 => x"fac21ec4",
  1582 => x"c149bfec",
  1583 => x"497487e1",
  1584 => x"87def7c0",
  1585 => x"c6e28ee4",
  1586 => x"1e731e87",
  1587 => x"fc494b71",
  1588 => x"497387d1",
  1589 => x"e187ccfc",
  1590 => x"731e87f9",
  1591 => x"c24b711e",
  1592 => x"d5024aa3",
  1593 => x"058ac187",
  1594 => x"fbc287db",
  1595 => x"d402bfc0",
  1596 => x"88c14887",
  1597 => x"58c4fbc2",
  1598 => x"fbc287cb",
  1599 => x"c148bfc0",
  1600 => x"c4fbc280",
  1601 => x"c01ec758",
  1602 => x"c4f7c11e",
  1603 => x"ecfac21e",
  1604 => x"87cb49bf",
  1605 => x"f6c04973",
  1606 => x"8ef487c8",
  1607 => x"0e87f4e0",
  1608 => x"5d5c5b5e",
  1609 => x"86d8ff0e",
  1610 => x"c859a6dc",
  1611 => x"78c048a6",
  1612 => x"78c080c4",
  1613 => x"c280c44d",
  1614 => x"78bfc0fb",
  1615 => x"c348d4ff",
  1616 => x"d0ff78ff",
  1617 => x"c0c848bf",
  1618 => x"a6c498c0",
  1619 => x"02987058",
  1620 => x"d0ff87d0",
  1621 => x"c0c848bf",
  1622 => x"a6c498c0",
  1623 => x"05987058",
  1624 => x"d0ff87f0",
  1625 => x"78e1c048",
  1626 => x"d448d4ff",
  1627 => x"d5ddff78",
  1628 => x"48d4ff87",
  1629 => x"d478ffc3",
  1630 => x"d4ff48a6",
  1631 => x"66d478bf",
  1632 => x"a8fbc048",
  1633 => x"87d3c102",
  1634 => x"4a66f8c0",
  1635 => x"7e6a82c4",
  1636 => x"d2c11e72",
  1637 => x"66c448d9",
  1638 => x"4aa1c849",
  1639 => x"aa714120",
  1640 => x"1087f905",
  1641 => x"c04a2651",
  1642 => x"c84966f8",
  1643 => x"f4dec181",
  1644 => x"c7496a79",
  1645 => x"5166d481",
  1646 => x"1ed81ec1",
  1647 => x"81c8496a",
  1648 => x"87d9dcff",
  1649 => x"66d086c8",
  1650 => x"a8b7c048",
  1651 => x"c187c401",
  1652 => x"d087c84d",
  1653 => x"88c14866",
  1654 => x"d458a6d4",
  1655 => x"f4ca0266",
  1656 => x"66c0c187",
  1657 => x"ca03adb7",
  1658 => x"d4ff87eb",
  1659 => x"78ffc348",
  1660 => x"ff48a6d4",
  1661 => x"d478bfd4",
  1662 => x"c6c14866",
  1663 => x"58a6c488",
  1664 => x"c0029870",
  1665 => x"c94887e6",
  1666 => x"58a6c488",
  1667 => x"c4029870",
  1668 => x"c14887d5",
  1669 => x"58a6c488",
  1670 => x"c1029870",
  1671 => x"c44887e3",
  1672 => x"7058a688",
  1673 => x"fec30298",
  1674 => x"87d3c987",
  1675 => x"c10566d8",
  1676 => x"d4ff87c5",
  1677 => x"78ffc348",
  1678 => x"1eca1ec0",
  1679 => x"93cc4b75",
  1680 => x"8366c0c1",
  1681 => x"6c4ca3c4",
  1682 => x"d0daff49",
  1683 => x"de1ec187",
  1684 => x"ff496c1e",
  1685 => x"d087c6da",
  1686 => x"49a3c886",
  1687 => x"79f4dec1",
  1688 => x"adb766d0",
  1689 => x"c187c504",
  1690 => x"87dac885",
  1691 => x"c14866d0",
  1692 => x"58a6d488",
  1693 => x"ff87cfc8",
  1694 => x"d887cbd9",
  1695 => x"c5c858a6",
  1696 => x"d2dbff87",
  1697 => x"58a6cc87",
  1698 => x"a8b766cc",
  1699 => x"cc87c606",
  1700 => x"66c848a6",
  1701 => x"fedaff78",
  1702 => x"a8ecc087",
  1703 => x"87c7c205",
  1704 => x"c10566d8",
  1705 => x"497587f7",
  1706 => x"f8c091cc",
  1707 => x"a1c48166",
  1708 => x"c14c6a4a",
  1709 => x"66c84aa1",
  1710 => x"7997c252",
  1711 => x"dfc181c8",
  1712 => x"d4ff79c2",
  1713 => x"78ffc348",
  1714 => x"ff48a6d4",
  1715 => x"d478bfd4",
  1716 => x"e8c00266",
  1717 => x"fbc04887",
  1718 => x"e0c002a8",
  1719 => x"9766d487",
  1720 => x"ff84c17c",
  1721 => x"ffc348d4",
  1722 => x"48a6d478",
  1723 => x"78bfd4ff",
  1724 => x"c80266d4",
  1725 => x"fbc04887",
  1726 => x"e0ff05a8",
  1727 => x"54e0c087",
  1728 => x"c054c1c2",
  1729 => x"66d07c97",
  1730 => x"c504adb7",
  1731 => x"c585c187",
  1732 => x"66d087f4",
  1733 => x"d488c148",
  1734 => x"e9c558a6",
  1735 => x"e5d6ff87",
  1736 => x"58a6d887",
  1737 => x"c887dfc5",
  1738 => x"66d84866",
  1739 => x"c4c505a8",
  1740 => x"48a6dc87",
  1741 => x"d8ff78c0",
  1742 => x"a6d887dd",
  1743 => x"d6d8ff58",
  1744 => x"a6e4c087",
  1745 => x"a8ecc058",
  1746 => x"87cac005",
  1747 => x"48a6e0c0",
  1748 => x"c07866d4",
  1749 => x"d4ff87c6",
  1750 => x"78ffc348",
  1751 => x"91cc4975",
  1752 => x"4866f8c0",
  1753 => x"a6c48071",
  1754 => x"c3496e58",
  1755 => x"5166d481",
  1756 => x"4966e0c0",
  1757 => x"66d481c1",
  1758 => x"7148c189",
  1759 => x"c1497030",
  1760 => x"c14a6e89",
  1761 => x"97097282",
  1762 => x"486e0979",
  1763 => x"fac250c2",
  1764 => x"d449bfe8",
  1765 => x"9729b766",
  1766 => x"71484a6a",
  1767 => x"a6e8c098",
  1768 => x"c4486e58",
  1769 => x"58a6c880",
  1770 => x"4cbf66c4",
  1771 => x"c84866d8",
  1772 => x"c002a866",
  1773 => x"e0c087c9",
  1774 => x"78c048a6",
  1775 => x"c087c6c0",
  1776 => x"c148a6e0",
  1777 => x"66e0c078",
  1778 => x"1ee0c01e",
  1779 => x"d4ff4974",
  1780 => x"86c887cb",
  1781 => x"c058a6d8",
  1782 => x"c106a8b7",
  1783 => x"66d487da",
  1784 => x"bf66c484",
  1785 => x"81e0c049",
  1786 => x"c14b8974",
  1787 => x"714ae2d2",
  1788 => x"87d7d7fe",
  1789 => x"66dc84c2",
  1790 => x"c080c148",
  1791 => x"c058a6e0",
  1792 => x"c14966e4",
  1793 => x"02a97081",
  1794 => x"c087c9c0",
  1795 => x"c048a6e0",
  1796 => x"87c6c078",
  1797 => x"48a6e0c0",
  1798 => x"e0c078c1",
  1799 => x"66c81e66",
  1800 => x"e0c049bf",
  1801 => x"71897481",
  1802 => x"ff49741e",
  1803 => x"c887eed2",
  1804 => x"a8b7c086",
  1805 => x"87fefe01",
  1806 => x"c00266dc",
  1807 => x"496e87d2",
  1808 => x"66dc81c2",
  1809 => x"c8496e51",
  1810 => x"e3dfc181",
  1811 => x"87cdc079",
  1812 => x"81c2496e",
  1813 => x"c8496e51",
  1814 => x"c9e3c181",
  1815 => x"b766d079",
  1816 => x"c5c004ad",
  1817 => x"c085c187",
  1818 => x"66d087dc",
  1819 => x"d488c148",
  1820 => x"d1c058a6",
  1821 => x"cdd1ff87",
  1822 => x"58a6d887",
  1823 => x"ff87c7c0",
  1824 => x"d887c3d1",
  1825 => x"66d458a6",
  1826 => x"87c9c002",
  1827 => x"b766c0c1",
  1828 => x"d5f504ad",
  1829 => x"adb7c787",
  1830 => x"87dcc003",
  1831 => x"91cc4975",
  1832 => x"8166f8c0",
  1833 => x"6a4aa1c4",
  1834 => x"c852c04a",
  1835 => x"c179c081",
  1836 => x"adb7c785",
  1837 => x"87e4ff04",
  1838 => x"c00266d8",
  1839 => x"f8c087eb",
  1840 => x"d4c14966",
  1841 => x"66f8c081",
  1842 => x"82d5c14a",
  1843 => x"51c252c0",
  1844 => x"4966f8c0",
  1845 => x"c181dcc1",
  1846 => x"c079c2df",
  1847 => x"c14966f8",
  1848 => x"d2c181d8",
  1849 => x"d6c079e5",
  1850 => x"66f8c087",
  1851 => x"81d8c149",
  1852 => x"79ecd2c1",
  1853 => x"4966f8c0",
  1854 => x"c281dcc1",
  1855 => x"c179cdde",
  1856 => x"c04adae3",
  1857 => x"c14966f8",
  1858 => x"797281e8",
  1859 => x"48bfd0ff",
  1860 => x"98c0c0c8",
  1861 => x"7058a6c4",
  1862 => x"d1c00298",
  1863 => x"bfd0ff87",
  1864 => x"c0c0c848",
  1865 => x"58a6c498",
  1866 => x"ff059870",
  1867 => x"d0ff87ef",
  1868 => x"78e0c048",
  1869 => x"ff4866cc",
  1870 => x"d0ff8ed8",
  1871 => x"c71e87d1",
  1872 => x"c11ec01e",
  1873 => x"c21ec4f7",
  1874 => x"49bfecfa",
  1875 => x"c187d0ef",
  1876 => x"c049c4f7",
  1877 => x"f487d6e8",
  1878 => x"1e4f268e",
  1879 => x"c287c6ca",
  1880 => x"c048c8fb",
  1881 => x"48d4ff50",
  1882 => x"c178ffc3",
  1883 => x"fe49f3d2",
  1884 => x"fe87f4d0",
  1885 => x"7087f0dd",
  1886 => x"87cd0298",
  1887 => x"87f0eafe",
  1888 => x"c4029870",
  1889 => x"c24ac187",
  1890 => x"724ac087",
  1891 => x"87c8029a",
  1892 => x"49c9d3c1",
  1893 => x"87cfd0fe",
  1894 => x"bfd8ecc2",
  1895 => x"c2d4ff49",
  1896 => x"c0fbc287",
  1897 => x"c278c048",
  1898 => x"c048ecfa",
  1899 => x"cdfe4978",
  1900 => x"87ddc387",
  1901 => x"c087c2c9",
  1902 => x"ff87e1e7",
  1903 => x"4f2687f6",
  1904 => x"000014d2",
  1905 => x"00000002",
  1906 => x"00002ed8",
  1907 => x"0000151f",
  1908 => x"00000002",
  1909 => x"00002ef6",
  1910 => x"0000151f",
  1911 => x"00000002",
  1912 => x"00002f14",
  1913 => x"0000151f",
  1914 => x"00000002",
  1915 => x"00002f32",
  1916 => x"0000151f",
  1917 => x"00000002",
  1918 => x"00002f50",
  1919 => x"0000151f",
  1920 => x"00000002",
  1921 => x"00002f6e",
  1922 => x"0000151f",
  1923 => x"00000002",
  1924 => x"00002f8c",
  1925 => x"0000151f",
  1926 => x"00000002",
  1927 => x"00000000",
  1928 => x"000017c2",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"000015b6",
  1932 => x"d5c11e1e",
  1933 => x"58a6c487",
  1934 => x"1e4f2626",
  1935 => x"f0fe4a71",
  1936 => x"cd78c048",
  1937 => x"c10a7a0a",
  1938 => x"fe49d1f9",
  1939 => x"2687d8cd",
  1940 => x"7465534f",
  1941 => x"6e616820",
  1942 => x"72656c64",
  1943 => x"6e49000a",
  1944 => x"746e6920",
  1945 => x"75727265",
  1946 => x"63207470",
  1947 => x"74736e6f",
  1948 => x"74637572",
  1949 => x"000a726f",
  1950 => x"def9c11e",
  1951 => x"e6ccfe49",
  1952 => x"f0f8c187",
  1953 => x"87f3fe49",
  1954 => x"fe1e4f26",
  1955 => x"2648bff0",
  1956 => x"f0fe1e4f",
  1957 => x"2678c148",
  1958 => x"f0fe1e4f",
  1959 => x"2678c048",
  1960 => x"4a711e4f",
  1961 => x"a2c47ac0",
  1962 => x"c879c049",
  1963 => x"79c049a2",
  1964 => x"c049a2cc",
  1965 => x"0e4f2679",
  1966 => x"0e5c5b5e",
  1967 => x"4c7186f8",
  1968 => x"cc49a4c8",
  1969 => x"486b4ba4",
  1970 => x"a6c480c1",
  1971 => x"c898cf58",
  1972 => x"486958a6",
  1973 => x"05a866c4",
  1974 => x"486b87d4",
  1975 => x"a6c480c1",
  1976 => x"c898cf58",
  1977 => x"486958a6",
  1978 => x"02a866c4",
  1979 => x"e8fe87ec",
  1980 => x"a4d0c187",
  1981 => x"c4486b49",
  1982 => x"58a6c490",
  1983 => x"66d48170",
  1984 => x"c1486b79",
  1985 => x"58a6c880",
  1986 => x"7b7098cf",
  1987 => x"fd87d2c1",
  1988 => x"8ef887ff",
  1989 => x"4d2687c2",
  1990 => x"4b264c26",
  1991 => x"5e0e4f26",
  1992 => x"0e5d5c5b",
  1993 => x"4d7186f8",
  1994 => x"6d4ca5c4",
  1995 => x"05a86c48",
  1996 => x"48ff87c5",
  1997 => x"fd87e5c0",
  1998 => x"a5d087df",
  1999 => x"c4486c4b",
  2000 => x"58a6c490",
  2001 => x"4b6b8370",
  2002 => x"6c9bffc3",
  2003 => x"c880c148",
  2004 => x"98cf58a6",
  2005 => x"f8fc7c70",
  2006 => x"48497387",
  2007 => x"f5fe8ef8",
  2008 => x"1e731e87",
  2009 => x"f0fc86f8",
  2010 => x"4bbfe087",
  2011 => x"c0e0c049",
  2012 => x"e7c00299",
  2013 => x"c34a7387",
  2014 => x"fec29aff",
  2015 => x"c448bfea",
  2016 => x"58a6c490",
  2017 => x"49fafec2",
  2018 => x"79728170",
  2019 => x"bfeafec2",
  2020 => x"c880c148",
  2021 => x"98cf58a6",
  2022 => x"58eefec2",
  2023 => x"c0d04973",
  2024 => x"f2c00299",
  2025 => x"f2fec287",
  2026 => x"fec248bf",
  2027 => x"02a8bff6",
  2028 => x"c287e4c0",
  2029 => x"48bff2fe",
  2030 => x"a6c490c4",
  2031 => x"faffc258",
  2032 => x"e0817049",
  2033 => x"c2786948",
  2034 => x"48bff2fe",
  2035 => x"a6c880c1",
  2036 => x"c298cf58",
  2037 => x"fa58f6fe",
  2038 => x"a6c487f0",
  2039 => x"87f1fa58",
  2040 => x"f5fc8ef8",
  2041 => x"fec21e87",
  2042 => x"f4fa49ea",
  2043 => x"e1fdc187",
  2044 => x"87c7f949",
  2045 => x"2687f5c3",
  2046 => x"1e731e4f",
  2047 => x"49eafec2",
  2048 => x"7087dbfc",
  2049 => x"aab7c04a",
  2050 => x"87ccc204",
  2051 => x"05aaf0c3",
  2052 => x"c2c287c9",
  2053 => x"78c148e4",
  2054 => x"c387edc1",
  2055 => x"c905aae0",
  2056 => x"e8c2c287",
  2057 => x"c178c148",
  2058 => x"c2c287de",
  2059 => x"c602bfe8",
  2060 => x"a2c0c287",
  2061 => x"7287c24b",
  2062 => x"e4c2c24b",
  2063 => x"e0c002bf",
  2064 => x"c4497387",
  2065 => x"c29129b7",
  2066 => x"7381ecc2",
  2067 => x"c29acf4a",
  2068 => x"7248c192",
  2069 => x"ff4a7030",
  2070 => x"694872ba",
  2071 => x"db797098",
  2072 => x"c4497387",
  2073 => x"c29129b7",
  2074 => x"7381ecc2",
  2075 => x"c29acf4a",
  2076 => x"7248c392",
  2077 => x"484a7030",
  2078 => x"7970b069",
  2079 => x"48e8c2c2",
  2080 => x"c2c278c0",
  2081 => x"78c048e4",
  2082 => x"49eafec2",
  2083 => x"7087cffa",
  2084 => x"aab7c04a",
  2085 => x"87f4fd03",
  2086 => x"87c448c0",
  2087 => x"4c264d26",
  2088 => x"4f264b26",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"724ac01e",
  2108 => x"c291c449",
  2109 => x"c081ecc2",
  2110 => x"d082c179",
  2111 => x"ee04aab7",
  2112 => x"0e4f2687",
  2113 => x"5d5c5b5e",
  2114 => x"f64d710e",
  2115 => x"4a7587cb",
  2116 => x"922ab7c4",
  2117 => x"82ecc2c2",
  2118 => x"9ccf4c75",
  2119 => x"496a94c2",
  2120 => x"c32b744b",
  2121 => x"7448c29b",
  2122 => x"ff4c7030",
  2123 => x"714874bc",
  2124 => x"f57a7098",
  2125 => x"487387db",
  2126 => x"1e87e1fd",
  2127 => x"bfd0ff1e",
  2128 => x"c0c0c848",
  2129 => x"58a6c498",
  2130 => x"d0029870",
  2131 => x"bfd0ff87",
  2132 => x"c0c0c848",
  2133 => x"58a6c498",
  2134 => x"f0059870",
  2135 => x"48d0ff87",
  2136 => x"7178e1c4",
  2137 => x"08d4ff48",
  2138 => x"4866c878",
  2139 => x"7808d4ff",
  2140 => x"1e4f2626",
  2141 => x"c84a711e",
  2142 => x"721e4966",
  2143 => x"87fbfe49",
  2144 => x"d0ff86c4",
  2145 => x"c0c848bf",
  2146 => x"a6c498c0",
  2147 => x"02987058",
  2148 => x"d0ff87d0",
  2149 => x"c0c848bf",
  2150 => x"a6c498c0",
  2151 => x"05987058",
  2152 => x"d0ff87f0",
  2153 => x"78e0c048",
  2154 => x"1e4f2626",
  2155 => x"4b711e73",
  2156 => x"731e66c8",
  2157 => x"a2e0c14a",
  2158 => x"87f7fe49",
  2159 => x"2687c426",
  2160 => x"264c264d",
  2161 => x"1e4f264b",
  2162 => x"bfd0ff1e",
  2163 => x"c0c0c848",
  2164 => x"58a6c498",
  2165 => x"d0029870",
  2166 => x"bfd0ff87",
  2167 => x"c0c0c848",
  2168 => x"58a6c498",
  2169 => x"f0059870",
  2170 => x"48d0ff87",
  2171 => x"7178c9c4",
  2172 => x"08d4ff48",
  2173 => x"4f262678",
  2174 => x"4a711e1e",
  2175 => x"87c7ff49",
  2176 => x"48bfd0ff",
  2177 => x"98c0c0c8",
  2178 => x"7058a6c4",
  2179 => x"87d00298",
  2180 => x"48bfd0ff",
  2181 => x"98c0c0c8",
  2182 => x"7058a6c4",
  2183 => x"87f00598",
  2184 => x"c848d0ff",
  2185 => x"4f262678",
  2186 => x"1e1e731e",
  2187 => x"c1c34b71",
  2188 => x"c302bfc6",
  2189 => x"87ccc387",
  2190 => x"48bfd0ff",
  2191 => x"98c0c0c8",
  2192 => x"7058a6c4",
  2193 => x"87d00298",
  2194 => x"48bfd0ff",
  2195 => x"98c0c0c8",
  2196 => x"7058a6c4",
  2197 => x"87f00598",
  2198 => x"c448d0ff",
  2199 => x"487378c9",
  2200 => x"ffb0e0c0",
  2201 => x"c37808d4",
  2202 => x"c048fac0",
  2203 => x"0266cc78",
  2204 => x"ffc387c5",
  2205 => x"c087c249",
  2206 => x"c2c1c349",
  2207 => x"0266d059",
  2208 => x"d5c587c6",
  2209 => x"87c44ad5",
  2210 => x"4affffcf",
  2211 => x"5ac6c1c3",
  2212 => x"48c6c1c3",
  2213 => x"c42678c1",
  2214 => x"264d2687",
  2215 => x"264b264c",
  2216 => x"5b5e0e4f",
  2217 => x"710e5d5c",
  2218 => x"c2c1c34a",
  2219 => x"9a724cbf",
  2220 => x"4987cb02",
  2221 => x"c9c291c8",
  2222 => x"83714be2",
  2223 => x"cdc287c4",
  2224 => x"4dc04be2",
  2225 => x"99744913",
  2226 => x"bffec0c3",
  2227 => x"ffb87148",
  2228 => x"c17808d4",
  2229 => x"c8852cb7",
  2230 => x"e704adb7",
  2231 => x"fac0c387",
  2232 => x"80c848bf",
  2233 => x"58fec0c3",
  2234 => x"1e87eefe",
  2235 => x"4b711e73",
  2236 => x"029a4a13",
  2237 => x"497287cb",
  2238 => x"1387e6fe",
  2239 => x"f5059a4a",
  2240 => x"87d9fe87",
  2241 => x"c0c31e1e",
  2242 => x"c349bffa",
  2243 => x"c148fac0",
  2244 => x"c0c478a1",
  2245 => x"db03a9b7",
  2246 => x"48d4ff87",
  2247 => x"bffec0c3",
  2248 => x"fac0c378",
  2249 => x"c0c349bf",
  2250 => x"a1c148fa",
  2251 => x"b7c0c478",
  2252 => x"87e504a9",
  2253 => x"48bfd0ff",
  2254 => x"98c0c0c8",
  2255 => x"7058a6c4",
  2256 => x"87d00298",
  2257 => x"48bfd0ff",
  2258 => x"98c0c0c8",
  2259 => x"7058a6c4",
  2260 => x"87f00598",
  2261 => x"c848d0ff",
  2262 => x"c6c1c378",
  2263 => x"2678c048",
  2264 => x"00004f26",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"005f5f00",
  2268 => x"03000000",
  2269 => x"03030003",
  2270 => x"7f140000",
  2271 => x"7f7f147f",
  2272 => x"24000014",
  2273 => x"3a6b6b2e",
  2274 => x"6a4c0012",
  2275 => x"566c1836",
  2276 => x"7e300032",
  2277 => x"3a77594f",
  2278 => x"00004068",
  2279 => x"00030704",
  2280 => x"00000000",
  2281 => x"41633e1c",
  2282 => x"00000000",
  2283 => x"1c3e6341",
  2284 => x"2a080000",
  2285 => x"3e1c1c3e",
  2286 => x"0800082a",
  2287 => x"083e3e08",
  2288 => x"00000008",
  2289 => x"0060e080",
  2290 => x"08000000",
  2291 => x"08080808",
  2292 => x"00000008",
  2293 => x"00606000",
  2294 => x"60400000",
  2295 => x"060c1830",
  2296 => x"3e000103",
  2297 => x"7f4d597f",
  2298 => x"0400003e",
  2299 => x"007f7f06",
  2300 => x"42000000",
  2301 => x"4f597163",
  2302 => x"22000046",
  2303 => x"7f494963",
  2304 => x"1c180036",
  2305 => x"7f7f1316",
  2306 => x"27000010",
  2307 => x"7d454567",
  2308 => x"3c000039",
  2309 => x"79494b7e",
  2310 => x"01000030",
  2311 => x"0f797101",
  2312 => x"36000007",
  2313 => x"7f49497f",
  2314 => x"06000036",
  2315 => x"3f69494f",
  2316 => x"0000001e",
  2317 => x"00666600",
  2318 => x"00000000",
  2319 => x"0066e680",
  2320 => x"08000000",
  2321 => x"22141408",
  2322 => x"14000022",
  2323 => x"14141414",
  2324 => x"22000014",
  2325 => x"08141422",
  2326 => x"02000008",
  2327 => x"0f595103",
  2328 => x"7f3e0006",
  2329 => x"1f555d41",
  2330 => x"7e00001e",
  2331 => x"7f09097f",
  2332 => x"7f00007e",
  2333 => x"7f49497f",
  2334 => x"1c000036",
  2335 => x"4141633e",
  2336 => x"7f000041",
  2337 => x"3e63417f",
  2338 => x"7f00001c",
  2339 => x"4149497f",
  2340 => x"7f000041",
  2341 => x"0109097f",
  2342 => x"3e000001",
  2343 => x"7b49417f",
  2344 => x"7f00007a",
  2345 => x"7f08087f",
  2346 => x"0000007f",
  2347 => x"417f7f41",
  2348 => x"20000000",
  2349 => x"7f404060",
  2350 => x"7f7f003f",
  2351 => x"63361c08",
  2352 => x"7f000041",
  2353 => x"4040407f",
  2354 => x"7f7f0040",
  2355 => x"7f060c06",
  2356 => x"7f7f007f",
  2357 => x"7f180c06",
  2358 => x"3e00007f",
  2359 => x"7f41417f",
  2360 => x"7f00003e",
  2361 => x"0f09097f",
  2362 => x"7f3e0006",
  2363 => x"7e7f6141",
  2364 => x"7f000040",
  2365 => x"7f19097f",
  2366 => x"26000066",
  2367 => x"7b594d6f",
  2368 => x"01000032",
  2369 => x"017f7f01",
  2370 => x"3f000001",
  2371 => x"7f40407f",
  2372 => x"0f00003f",
  2373 => x"3f70703f",
  2374 => x"7f7f000f",
  2375 => x"7f301830",
  2376 => x"6341007f",
  2377 => x"361c1c36",
  2378 => x"03014163",
  2379 => x"067c7c06",
  2380 => x"71610103",
  2381 => x"43474d59",
  2382 => x"00000041",
  2383 => x"41417f7f",
  2384 => x"03010000",
  2385 => x"30180c06",
  2386 => x"00004060",
  2387 => x"7f7f4141",
  2388 => x"0c080000",
  2389 => x"0c060306",
  2390 => x"80800008",
  2391 => x"80808080",
  2392 => x"00000080",
  2393 => x"04070300",
  2394 => x"20000000",
  2395 => x"7c545474",
  2396 => x"7f000078",
  2397 => x"7c44447f",
  2398 => x"38000038",
  2399 => x"4444447c",
  2400 => x"38000000",
  2401 => x"7f44447c",
  2402 => x"3800007f",
  2403 => x"5c54547c",
  2404 => x"04000018",
  2405 => x"05057f7e",
  2406 => x"18000000",
  2407 => x"fca4a4bc",
  2408 => x"7f00007c",
  2409 => x"7c04047f",
  2410 => x"00000078",
  2411 => x"407d3d00",
  2412 => x"80000000",
  2413 => x"7dfd8080",
  2414 => x"7f000000",
  2415 => x"6c38107f",
  2416 => x"00000044",
  2417 => x"407f3f00",
  2418 => x"7c7c0000",
  2419 => x"7c0c180c",
  2420 => x"7c000078",
  2421 => x"7c04047c",
  2422 => x"38000078",
  2423 => x"7c44447c",
  2424 => x"fc000038",
  2425 => x"3c2424fc",
  2426 => x"18000018",
  2427 => x"fc24243c",
  2428 => x"7c0000fc",
  2429 => x"0c04047c",
  2430 => x"48000008",
  2431 => x"7454545c",
  2432 => x"04000020",
  2433 => x"44447f3f",
  2434 => x"3c000000",
  2435 => x"7c40407c",
  2436 => x"1c00007c",
  2437 => x"3c60603c",
  2438 => x"7c3c001c",
  2439 => x"7c603060",
  2440 => x"6c44003c",
  2441 => x"6c381038",
  2442 => x"1c000044",
  2443 => x"3c60e0bc",
  2444 => x"4400001c",
  2445 => x"4c5c7464",
  2446 => x"08000044",
  2447 => x"41773e08",
  2448 => x"00000041",
  2449 => x"007f7f00",
  2450 => x"41000000",
  2451 => x"083e7741",
  2452 => x"01020008",
  2453 => x"02020301",
  2454 => x"7f7f0001",
  2455 => x"7f7f7f7f",
  2456 => x"0808007f",
  2457 => x"3e3e1c1c",
  2458 => x"7f7f7f7f",
  2459 => x"1c1c3e3e",
  2460 => x"10000808",
  2461 => x"187c7c18",
  2462 => x"10000010",
  2463 => x"307c7c30",
  2464 => x"30100010",
  2465 => x"1e786060",
  2466 => x"66420006",
  2467 => x"663c183c",
  2468 => x"38780042",
  2469 => x"6cc6c26a",
  2470 => x"00600038",
  2471 => x"00006000",
  2472 => x"5e0e0060",
  2473 => x"0e5d5c5b",
  2474 => x"c34c711e",
  2475 => x"4bbfcec1",
  2476 => x"48d2c1c3",
  2477 => x"1e7478c0",
  2478 => x"1efddcc2",
  2479 => x"87fce6fd",
  2480 => x"6b9786c8",
  2481 => x"c1029949",
  2482 => x"1ec087c6",
  2483 => x"c348a6c4",
  2484 => x"78bfd2c1",
  2485 => x"02ac66c4",
  2486 => x"4dc087c4",
  2487 => x"4dc187c2",
  2488 => x"66c81e75",
  2489 => x"87c0ed49",
  2490 => x"e0c086c8",
  2491 => x"87f1ee49",
  2492 => x"6a4aa3c4",
  2493 => x"87f3ef49",
  2494 => x"c387c9f0",
  2495 => x"48bfd2c1",
  2496 => x"c1c380c1",
  2497 => x"83cc58d6",
  2498 => x"99496b97",
  2499 => x"87fafe05",
  2500 => x"bfd2c1c3",
  2501 => x"adb7c84d",
  2502 => x"c087d903",
  2503 => x"c1c31e1e",
  2504 => x"ec49bfd2",
  2505 => x"86c887c2",
  2506 => x"c187d9ef",
  2507 => x"adb7c885",
  2508 => x"87e7ff04",
  2509 => x"264d2626",
  2510 => x"264b264c",
  2511 => x"6769484f",
  2512 => x"67696c68",
  2513 => x"72207468",
  2514 => x"2520776f",
  2515 => x"4d000a64",
  2516 => x"20756e65",
  2517 => x"69736976",
  2518 => x"20656c62",
  2519 => x"000a6425",
  2520 => x"6c6c6143",
  2521 => x"6b636162",
  2522 => x"0a782520",
  2523 => x"4a711e00",
  2524 => x"5ad2c1c3",
  2525 => x"bfd6c1c3",
  2526 => x"87e6fc49",
  2527 => x"bfd2c1c3",
  2528 => x"c389c149",
  2529 => x"7159dac1",
  2530 => x"2687d7fc",
  2531 => x"c0c11e4f",
  2532 => x"87e4e949",
  2533 => x"48c1ecc2",
  2534 => x"4f2678c0",
  2535 => x"5c5b5e0e",
  2536 => x"86f40e5d",
  2537 => x"c048a6c8",
  2538 => x"7ebfec78",
  2539 => x"c1c380fc",
  2540 => x"c378bfce",
  2541 => x"4dbfdac1",
  2542 => x"c74cbfe8",
  2543 => x"87c3e549",
  2544 => x"99c24970",
  2545 => x"c287cf05",
  2546 => x"49bff9eb",
  2547 => x"996eb9ff",
  2548 => x"c00299c1",
  2549 => x"49c787fd",
  2550 => x"7087e8e4",
  2551 => x"87cd0298",
  2552 => x"c787d6e0",
  2553 => x"87dbe449",
  2554 => x"f3059870",
  2555 => x"c1ecc287",
  2556 => x"ddc21ebf",
  2557 => x"e2fd1ecf",
  2558 => x"86c887c2",
  2559 => x"bfc1ecc2",
  2560 => x"c2bac14a",
  2561 => x"c15ac5ec",
  2562 => x"e749a2c0",
  2563 => x"a6c887ea",
  2564 => x"c278c148",
  2565 => x"6e48f9eb",
  2566 => x"c1ecc278",
  2567 => x"dac105bf",
  2568 => x"48a6c487",
  2569 => x"78c0c0c8",
  2570 => x"7ec5ecc2",
  2571 => x"49bf976e",
  2572 => x"80c1486e",
  2573 => x"7158a6c4",
  2574 => x"7087c8e3",
  2575 => x"87c30298",
  2576 => x"c4b466c4",
  2577 => x"b7c14866",
  2578 => x"58a6c828",
  2579 => x"ff059870",
  2580 => x"497487da",
  2581 => x"7199ffc3",
  2582 => x"e549c01e",
  2583 => x"497487cd",
  2584 => x"7129b7c8",
  2585 => x"e549c11e",
  2586 => x"86c887c1",
  2587 => x"e249fdc3",
  2588 => x"fac387d1",
  2589 => x"87cbe249",
  2590 => x"7487e9c9",
  2591 => x"99ffc349",
  2592 => x"712cb7c8",
  2593 => x"029c74b4",
  2594 => x"c8ff87df",
  2595 => x"496e7ebf",
  2596 => x"bffdebc2",
  2597 => x"a9c0c289",
  2598 => x"87c4c003",
  2599 => x"87cf4cc0",
  2600 => x"48fdebc2",
  2601 => x"c6c0786e",
  2602 => x"fdebc287",
  2603 => x"7478c048",
  2604 => x"0599c849",
  2605 => x"f5c387ce",
  2606 => x"87c7e149",
  2607 => x"99c24970",
  2608 => x"87eec002",
  2609 => x"bfd6c1c3",
  2610 => x"87c9c002",
  2611 => x"c388c148",
  2612 => x"d858dac1",
  2613 => x"d2c1c387",
  2614 => x"91cc49bf",
  2615 => x"c88166c4",
  2616 => x"bf6e7ea1",
  2617 => x"87c5c002",
  2618 => x"7349ff4b",
  2619 => x"48a6c80f",
  2620 => x"497478c1",
  2621 => x"c00599c4",
  2622 => x"f2c387ce",
  2623 => x"87c3e049",
  2624 => x"99c24970",
  2625 => x"87fec002",
  2626 => x"c348a6c8",
  2627 => x"78bfd2c1",
  2628 => x"c14966c8",
  2629 => x"d6c1c389",
  2630 => x"b76e7ebf",
  2631 => x"cac006a9",
  2632 => x"80c14887",
  2633 => x"58dac1c3",
  2634 => x"c887d6c0",
  2635 => x"91cc4966",
  2636 => x"c88166c4",
  2637 => x"bf6e7ea1",
  2638 => x"87c5c002",
  2639 => x"7349fe4b",
  2640 => x"48a6c80f",
  2641 => x"fdc378c1",
  2642 => x"f6deff49",
  2643 => x"c2497087",
  2644 => x"eec00299",
  2645 => x"d6c1c387",
  2646 => x"c9c002bf",
  2647 => x"d6c1c387",
  2648 => x"c078c048",
  2649 => x"c1c387d8",
  2650 => x"cc49bfd2",
  2651 => x"8166c491",
  2652 => x"6e7ea1c8",
  2653 => x"c5c002bf",
  2654 => x"49fd4b87",
  2655 => x"a6c80f73",
  2656 => x"c378c148",
  2657 => x"ddff49fa",
  2658 => x"497087f9",
  2659 => x"c10299c2",
  2660 => x"a6c887c0",
  2661 => x"d2c1c348",
  2662 => x"66c878bf",
  2663 => x"c488c148",
  2664 => x"c1c358a6",
  2665 => x"6e48bfd6",
  2666 => x"c003a8b7",
  2667 => x"c1c387c9",
  2668 => x"786e48d6",
  2669 => x"c887d6c0",
  2670 => x"91cc4966",
  2671 => x"c88166c4",
  2672 => x"bf6e7ea1",
  2673 => x"87c5c002",
  2674 => x"7349fc4b",
  2675 => x"48a6c80f",
  2676 => x"c1c378c1",
  2677 => x"c04bbfd6",
  2678 => x"c006abb7",
  2679 => x"8bc187c9",
  2680 => x"01abb7c0",
  2681 => x"7487f7ff",
  2682 => x"99f0c349",
  2683 => x"87cfc005",
  2684 => x"ff49dac1",
  2685 => x"7087ccdc",
  2686 => x"0299c249",
  2687 => x"c387e8c2",
  2688 => x"7ebfcec1",
  2689 => x"bfd6c1c3",
  2690 => x"abb7c04b",
  2691 => x"87d0c006",
  2692 => x"80cc486e",
  2693 => x"c158a6c4",
  2694 => x"abb7c08b",
  2695 => x"87f0ff01",
  2696 => x"4abf976e",
  2697 => x"c0028ac1",
  2698 => x"028a87f7",
  2699 => x"8a87d6c0",
  2700 => x"87cac102",
  2701 => x"eec1058a",
  2702 => x"c84a6e87",
  2703 => x"f4496a82",
  2704 => x"e2c187eb",
  2705 => x"c84b6e87",
  2706 => x"c21e6b83",
  2707 => x"fd1ee0dd",
  2708 => x"c887e9d8",
  2709 => x"c34b6b86",
  2710 => x"49bfd6c1",
  2711 => x"c6c10f73",
  2712 => x"c8496e87",
  2713 => x"6948c181",
  2714 => x"c3497030",
  2715 => x"48bfcac1",
  2716 => x"c1c3b871",
  2717 => x"a6c858ce",
  2718 => x"c078c148",
  2719 => x"496e87e9",
  2720 => x"486e81c8",
  2721 => x"a6c880cb",
  2722 => x"9766c458",
  2723 => x"a2c14abf",
  2724 => x"4969974b",
  2725 => x"c004abb7",
  2726 => x"4bc087c2",
  2727 => x"970b66c4",
  2728 => x"a6c80b7b",
  2729 => x"7578c148",
  2730 => x"e9c0029d",
  2731 => x"c0026d87",
  2732 => x"496d87e4",
  2733 => x"87cbd9ff",
  2734 => x"99c14970",
  2735 => x"87cbc002",
  2736 => x"c34ba5c4",
  2737 => x"49bfd6c1",
  2738 => x"c80f4b6b",
  2739 => x"c5c00285",
  2740 => x"ff056d87",
  2741 => x"66c887dc",
  2742 => x"87c8c002",
  2743 => x"bfd6c1c3",
  2744 => x"87feee49",
  2745 => x"ccf18ef4",
  2746 => x"11125887",
  2747 => x"1c1b1d14",
  2748 => x"91595a23",
  2749 => x"ebf2f594",
  2750 => x"000000f4",
  2751 => x"00000000",
  2752 => x"00000000",
  2753 => x"14125800",
  2754 => x"1c1b1d11",
  2755 => x"94595a23",
  2756 => x"ebf2f591",
  2757 => x"000000f4",
  2758 => x"00002b1c",
  2759 => x"4f545541",
  2760 => x"544f4f42",
  2761 => x"0053454e",
  2762 => x"00001e78",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
