library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c8ecc287",
    12 => x"86c0c44e",
    13 => x"49c8ecc2",
    14 => x"48d4d7c2",
    15 => x"0389d089",
    16 => x"404040c0",
    17 => x"d087f640",
    18 => x"50c00581",
    19 => x"f90589c1",
    20 => x"d4d7c287",
    21 => x"d0d7c24d",
    22 => x"02ad744c",
    23 => x"0f2487c4",
    24 => x"e1c187f7",
    25 => x"d7c287c1",
    26 => x"d7c24dd4",
    27 => x"ad744cd4",
    28 => x"c487c602",
    29 => x"f50f6c8c",
    30 => x"87fd0087",
    31 => x"5c5b5e0e",
    32 => x"c04b710e",
    33 => x"9a4a134c",
    34 => x"7287cd02",
    35 => x"87e0c049",
    36 => x"4a1384c1",
    37 => x"87f3059a",
    38 => x"4c264874",
    39 => x"4f264b26",
    40 => x"8148731e",
    41 => x"c502a973",
    42 => x"05531287",
    43 => x"4f2687f6",
    44 => x"c0ff1e1e",
    45 => x"c4486a4a",
    46 => x"a6c498c0",
    47 => x"02987058",
    48 => x"7a7187f3",
    49 => x"4f262648",
    50 => x"ff1e731e",
    51 => x"ffc34bd4",
    52 => x"c34a6b7b",
    53 => x"496b7bff",
    54 => x"b17232c8",
    55 => x"6b7bffc3",
    56 => x"7131c84a",
    57 => x"7bffc3b2",
    58 => x"32c8496b",
    59 => x"4871b172",
    60 => x"4d2687c4",
    61 => x"4b264c26",
    62 => x"5e0e4f26",
    63 => x"0e5d5c5b",
    64 => x"d4ff4a71",
    65 => x"c348724c",
    66 => x"7c7098ff",
    67 => x"bfd4d7c2",
    68 => x"d087c805",
    69 => x"30c94866",
    70 => x"d058a6d4",
    71 => x"29d84966",
    72 => x"ffc34871",
    73 => x"d07c7098",
    74 => x"29d04966",
    75 => x"ffc34871",
    76 => x"d07c7098",
    77 => x"29c84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"ffc34866",
    81 => x"727c7098",
    82 => x"7129d049",
    83 => x"98ffc348",
    84 => x"4b6c7c70",
    85 => x"4dfff0c9",
    86 => x"05abffc3",
    87 => x"ffc387d0",
    88 => x"c14b6c7c",
    89 => x"87c6028d",
    90 => x"02abffc3",
    91 => x"487387f0",
    92 => x"1e87fffd",
    93 => x"d4ff49c0",
    94 => x"78ffc348",
    95 => x"c8c381c1",
    96 => x"f104a9b7",
    97 => x"1e4f2687",
    98 => x"87e71e73",
    99 => x"4bdff8c4",
   100 => x"ffc01ec0",
   101 => x"49f7c1f0",
   102 => x"c487dffd",
   103 => x"05a8c186",
   104 => x"ff87eac0",
   105 => x"ffc348d4",
   106 => x"c0c0c178",
   107 => x"1ec0c0c0",
   108 => x"c1f0e1c0",
   109 => x"c1fd49e9",
   110 => x"7086c487",
   111 => x"87ca0598",
   112 => x"c348d4ff",
   113 => x"48c178ff",
   114 => x"e6fe87cb",
   115 => x"058bc187",
   116 => x"c087fdfe",
   117 => x"87defc48",
   118 => x"ff1e731e",
   119 => x"ffc348d4",
   120 => x"49d3c878",
   121 => x"d387d5fa",
   122 => x"c01ec04b",
   123 => x"c1c1f0ff",
   124 => x"87c6fc49",
   125 => x"987086c4",
   126 => x"ff87ca05",
   127 => x"ffc348d4",
   128 => x"cb48c178",
   129 => x"87ebfd87",
   130 => x"ff058bc1",
   131 => x"48c087db",
   132 => x"4387e3fb",
   133 => x"5300444d",
   134 => x"20434844",
   135 => x"6c696166",
   136 => x"49000a21",
   137 => x"00525245",
   138 => x"00495053",
   139 => x"74697257",
   140 => x"61662065",
   141 => x"64656c69",
   142 => x"5e0e000a",
   143 => x"ff0e5c5b",
   144 => x"eefc4cd4",
   145 => x"1eeac687",
   146 => x"c1f0e1c0",
   147 => x"e9fa49c8",
   148 => x"c186c487",
   149 => x"87c802a8",
   150 => x"c087fdfd",
   151 => x"87e8c148",
   152 => x"7087e5f9",
   153 => x"ffffcf49",
   154 => x"a9eac699",
   155 => x"fd87c802",
   156 => x"48c087e6",
   157 => x"c387d1c1",
   158 => x"f1c07cff",
   159 => x"87c7fc4b",
   160 => x"c0029870",
   161 => x"1ec087eb",
   162 => x"c1f0ffc0",
   163 => x"e9f949fa",
   164 => x"7086c487",
   165 => x"87d90598",
   166 => x"6c7cffc3",
   167 => x"7cffc349",
   168 => x"c17c7c7c",
   169 => x"c40299c0",
   170 => x"db48c187",
   171 => x"d748c087",
   172 => x"05abc287",
   173 => x"d7c887ca",
   174 => x"87c0f749",
   175 => x"87c848c0",
   176 => x"fe058bc1",
   177 => x"48c087f7",
   178 => x"0e87e9f8",
   179 => x"5d5c5b5e",
   180 => x"d0ff1e0e",
   181 => x"c0c0c84d",
   182 => x"d4d7c24b",
   183 => x"c878c148",
   184 => x"d7f649e8",
   185 => x"6d4cc787",
   186 => x"c4987348",
   187 => x"987058a6",
   188 => x"6d87cc02",
   189 => x"c4987348",
   190 => x"987058a6",
   191 => x"c287f405",
   192 => x"87eff97d",
   193 => x"9873486d",
   194 => x"7058a6c4",
   195 => x"87cc0298",
   196 => x"9873486d",
   197 => x"7058a6c4",
   198 => x"87f40598",
   199 => x"1ec07dc3",
   200 => x"c1d0e5c0",
   201 => x"d1f749c0",
   202 => x"c186c487",
   203 => x"87c105a8",
   204 => x"05acc24c",
   205 => x"e3c887cb",
   206 => x"87c0f549",
   207 => x"cec148c0",
   208 => x"058cc187",
   209 => x"fb87e0fe",
   210 => x"d7c287f0",
   211 => x"987058d8",
   212 => x"c187cd05",
   213 => x"f0ffc01e",
   214 => x"f649d0c1",
   215 => x"86c487dc",
   216 => x"c348d4ff",
   217 => x"ddc578ff",
   218 => x"dcd7c287",
   219 => x"73486d58",
   220 => x"58a6c498",
   221 => x"cc029870",
   222 => x"73486d87",
   223 => x"58a6c498",
   224 => x"f4059870",
   225 => x"ff7dc287",
   226 => x"ffc348d4",
   227 => x"2648c178",
   228 => x"0e87dff5",
   229 => x"5d5c5b5e",
   230 => x"c0c81e0e",
   231 => x"4cc04bc0",
   232 => x"dfcdeec5",
   233 => x"5ca6c44a",
   234 => x"c34cd4ff",
   235 => x"486c7cff",
   236 => x"05a8fec3",
   237 => x"7187c0c2",
   238 => x"e2c00599",
   239 => x"bfd0ff87",
   240 => x"c4987348",
   241 => x"987058a6",
   242 => x"ff87ce02",
   243 => x"7348bfd0",
   244 => x"58a6c498",
   245 => x"f2059870",
   246 => x"48d0ff87",
   247 => x"d478d1c4",
   248 => x"b7c04866",
   249 => x"e0c006a8",
   250 => x"7cffc387",
   251 => x"99714a6c",
   252 => x"7187c702",
   253 => x"0a7a970a",
   254 => x"66d481c1",
   255 => x"d888c148",
   256 => x"b7c058a6",
   257 => x"e0ff01a8",
   258 => x"7cffc387",
   259 => x"0599717c",
   260 => x"ff87e1c0",
   261 => x"7348bfd0",
   262 => x"58a6c498",
   263 => x"ce029870",
   264 => x"bfd0ff87",
   265 => x"c4987348",
   266 => x"987058a6",
   267 => x"ff87f205",
   268 => x"78d048d0",
   269 => x"c17e4ac1",
   270 => x"eefd058a",
   271 => x"26486e87",
   272 => x"0e87eff2",
   273 => x"0e5c5b5e",
   274 => x"c84a711e",
   275 => x"c04bc0c0",
   276 => x"48d4ff4c",
   277 => x"ff78ffc3",
   278 => x"7348bfd0",
   279 => x"58a6c498",
   280 => x"ce029870",
   281 => x"bfd0ff87",
   282 => x"c4987348",
   283 => x"987058a6",
   284 => x"ff87f205",
   285 => x"c3c448d0",
   286 => x"48d4ff78",
   287 => x"7278ffc3",
   288 => x"f0ffc01e",
   289 => x"f149d1c1",
   290 => x"86c487f0",
   291 => x"c0059870",
   292 => x"c0c887ee",
   293 => x"4966d41e",
   294 => x"c487f8fb",
   295 => x"ff4c7086",
   296 => x"7348bfd0",
   297 => x"58a6c498",
   298 => x"ce029870",
   299 => x"bfd0ff87",
   300 => x"c4987348",
   301 => x"987058a6",
   302 => x"ff87f205",
   303 => x"78c248d0",
   304 => x"f0264874",
   305 => x"5e0e87ee",
   306 => x"0e5d5c5b",
   307 => x"ffc01ec0",
   308 => x"49c9c1f0",
   309 => x"d287e3f0",
   310 => x"e2d7c21e",
   311 => x"87f3fa49",
   312 => x"4cc086c8",
   313 => x"b7d284c1",
   314 => x"87f804ac",
   315 => x"97e2d7c2",
   316 => x"c0c349bf",
   317 => x"a9c0c199",
   318 => x"87e7c005",
   319 => x"97e9d7c2",
   320 => x"31d049bf",
   321 => x"97ead7c2",
   322 => x"32c84abf",
   323 => x"d7c2b172",
   324 => x"4abf97eb",
   325 => x"cf4c71b1",
   326 => x"9cffffff",
   327 => x"34ca84c1",
   328 => x"c287e7c1",
   329 => x"bf97ebd7",
   330 => x"c631c149",
   331 => x"ecd7c299",
   332 => x"c74abf97",
   333 => x"b1722ab7",
   334 => x"97e7d7c2",
   335 => x"cf4d4abf",
   336 => x"e8d7c29d",
   337 => x"c34abf97",
   338 => x"c232ca9a",
   339 => x"bf97e9d7",
   340 => x"7333c24b",
   341 => x"ead7c2b2",
   342 => x"c34bbf97",
   343 => x"b7c69bc0",
   344 => x"c2b2732b",
   345 => x"7148c181",
   346 => x"c1497030",
   347 => x"70307548",
   348 => x"c14c724d",
   349 => x"c8947184",
   350 => x"06adb7c0",
   351 => x"34c187cc",
   352 => x"c0c82db7",
   353 => x"ff01adb7",
   354 => x"487487f4",
   355 => x"0e87e3ed",
   356 => x"0e5c5b5e",
   357 => x"4cc04b71",
   358 => x"c04866d0",
   359 => x"c006a8b7",
   360 => x"4a1387e3",
   361 => x"bf9766cc",
   362 => x"4866cc49",
   363 => x"a6d080c1",
   364 => x"aab77158",
   365 => x"c187c402",
   366 => x"c187cc48",
   367 => x"b766d084",
   368 => x"ddff04ac",
   369 => x"c248c087",
   370 => x"264d2687",
   371 => x"264b264c",
   372 => x"5b5e0e4f",
   373 => x"c20e5d5c",
   374 => x"c048c8e0",
   375 => x"c0d8c278",
   376 => x"f949c01e",
   377 => x"86c487dd",
   378 => x"c5059870",
   379 => x"c848c087",
   380 => x"4bc087ef",
   381 => x"48c0e5c2",
   382 => x"1ec878c1",
   383 => x"1eede0c0",
   384 => x"49f6d8c2",
   385 => x"c887c8fe",
   386 => x"05987086",
   387 => x"e5c287c6",
   388 => x"78c048c0",
   389 => x"e0c01ec8",
   390 => x"d9c21ef6",
   391 => x"eefd49d2",
   392 => x"7086c887",
   393 => x"87c60598",
   394 => x"48c0e5c2",
   395 => x"e5c278c0",
   396 => x"c002bfc0",
   397 => x"dfc287fa",
   398 => x"c24bbfc6",
   399 => x"bf9ffedf",
   400 => x"ead6c54a",
   401 => x"87c705aa",
   402 => x"bfc6dfc2",
   403 => x"ca87cc4b",
   404 => x"02aad5e9",
   405 => x"48c087c5",
   406 => x"c287c6c7",
   407 => x"731ec0d8",
   408 => x"87dff749",
   409 => x"987086c4",
   410 => x"c087c505",
   411 => x"87f1c648",
   412 => x"e0c01ec8",
   413 => x"d9c21eff",
   414 => x"d2fc49d2",
   415 => x"7086c887",
   416 => x"87c80598",
   417 => x"48c8e0c2",
   418 => x"87da78c1",
   419 => x"e1c01ec8",
   420 => x"d8c21ec8",
   421 => x"f6fb49f6",
   422 => x"7086c887",
   423 => x"c5c00298",
   424 => x"c548c087",
   425 => x"dfc287fb",
   426 => x"49bf97fe",
   427 => x"05a9d5c1",
   428 => x"c287cdc0",
   429 => x"bf97ffdf",
   430 => x"a9eac249",
   431 => x"87c5c002",
   432 => x"dcc548c0",
   433 => x"c0d8c287",
   434 => x"c34cbf97",
   435 => x"c002ace9",
   436 => x"ebc387cc",
   437 => x"c5c002ac",
   438 => x"c548c087",
   439 => x"d8c287c3",
   440 => x"49bf97cb",
   441 => x"ccc00599",
   442 => x"ccd8c287",
   443 => x"c249bf97",
   444 => x"c5c002a9",
   445 => x"c448c087",
   446 => x"d8c287e7",
   447 => x"48bf97cd",
   448 => x"58c4e0c2",
   449 => x"e0c288c1",
   450 => x"d8c258c8",
   451 => x"49bf97ce",
   452 => x"d8c28173",
   453 => x"4abf97cf",
   454 => x"7135c84d",
   455 => x"e0e4c285",
   456 => x"d0d8c25d",
   457 => x"c248bf97",
   458 => x"c258f4e4",
   459 => x"02bfc8e0",
   460 => x"c887dcc2",
   461 => x"e4e0c01e",
   462 => x"d2d9c21e",
   463 => x"87cff949",
   464 => x"987086c8",
   465 => x"87c5c002",
   466 => x"d4c348c0",
   467 => x"c0e0c287",
   468 => x"c4484abf",
   469 => x"d0e0c230",
   470 => x"f0e4c258",
   471 => x"e5d8c25a",
   472 => x"c849bf97",
   473 => x"e4d8c231",
   474 => x"a14bbf97",
   475 => x"e6d8c249",
   476 => x"d04bbf97",
   477 => x"49a17333",
   478 => x"97e7d8c2",
   479 => x"33d84bbf",
   480 => x"c249a173",
   481 => x"c259f8e4",
   482 => x"91bff0e4",
   483 => x"bfdce4c2",
   484 => x"e4e4c281",
   485 => x"edd8c259",
   486 => x"c84bbf97",
   487 => x"ecd8c233",
   488 => x"a34cbf97",
   489 => x"eed8c24b",
   490 => x"d04cbf97",
   491 => x"4ba37434",
   492 => x"97efd8c2",
   493 => x"9ccf4cbf",
   494 => x"a37434d8",
   495 => x"e8e4c24b",
   496 => x"738bc25b",
   497 => x"e8e4c292",
   498 => x"78a17248",
   499 => x"c287cbc1",
   500 => x"bf97d2d8",
   501 => x"c231c849",
   502 => x"bf97d1d8",
   503 => x"c249a14a",
   504 => x"c559d0e0",
   505 => x"81ffc731",
   506 => x"e4c229c9",
   507 => x"d8c259f0",
   508 => x"4abf97d7",
   509 => x"d8c232c8",
   510 => x"4bbf97d6",
   511 => x"e4c24aa2",
   512 => x"e4c25af8",
   513 => x"7592bff0",
   514 => x"ece4c282",
   515 => x"e4e4c25a",
   516 => x"c278c048",
   517 => x"7248e0e4",
   518 => x"49c078a1",
   519 => x"c187f7c7",
   520 => x"87e5f648",
   521 => x"33544146",
   522 => x"20202032",
   523 => x"54414600",
   524 => x"20203631",
   525 => x"41460020",
   526 => x"20323354",
   527 => x"46002020",
   528 => x"32335441",
   529 => x"00202020",
   530 => x"31544146",
   531 => x"20202036",
   532 => x"5b5e0e00",
   533 => x"710e5d5c",
   534 => x"c8e0c24a",
   535 => x"87cc02bf",
   536 => x"b7c74b72",
   537 => x"c14d722b",
   538 => x"87ca9dff",
   539 => x"b7c84b72",
   540 => x"c34d722b",
   541 => x"d8c29dff",
   542 => x"e4c21ec0",
   543 => x"7349bfdc",
   544 => x"feee7181",
   545 => x"7086c487",
   546 => x"87c50598",
   547 => x"e6c048c0",
   548 => x"c8e0c287",
   549 => x"87d202bf",
   550 => x"91c44975",
   551 => x"81c0d8c2",
   552 => x"ffcf4c69",
   553 => x"9cffffff",
   554 => x"497587cb",
   555 => x"d8c291c2",
   556 => x"699f81c0",
   557 => x"f448744c",
   558 => x"5e0e87cf",
   559 => x"0e5d5c5b",
   560 => x"4c7186f4",
   561 => x"e4c24bc0",
   562 => x"c47ebff8",
   563 => x"e4c248a6",
   564 => x"c878bffc",
   565 => x"78c048a6",
   566 => x"bfcce0c2",
   567 => x"06a8c048",
   568 => x"c887ddc2",
   569 => x"99cf4966",
   570 => x"c287d805",
   571 => x"c81ec0d8",
   572 => x"c1484966",
   573 => x"58a6cc80",
   574 => x"c487c8ed",
   575 => x"c0d8c286",
   576 => x"c087c34b",
   577 => x"6b9783e0",
   578 => x"c1029a4a",
   579 => x"e5c387e1",
   580 => x"dac102aa",
   581 => x"49a3cb87",
   582 => x"d8496997",
   583 => x"cec10599",
   584 => x"c01ecb87",
   585 => x"731e66e0",
   586 => x"87e3f149",
   587 => x"987086c8",
   588 => x"87fbc005",
   589 => x"c44aa3dc",
   590 => x"796a49a4",
   591 => x"c849a3da",
   592 => x"699f4da4",
   593 => x"e0c27d48",
   594 => x"d302bfc8",
   595 => x"49a3d487",
   596 => x"c049699f",
   597 => x"7199ffff",
   598 => x"c430d048",
   599 => x"87c258a6",
   600 => x"486e7ec0",
   601 => x"7d70806d",
   602 => x"48c17cc0",
   603 => x"c887c5c1",
   604 => x"80c14866",
   605 => x"c258a6cc",
   606 => x"a8bfcce0",
   607 => x"87e3fd04",
   608 => x"bfc8e0c2",
   609 => x"87eac002",
   610 => x"c4fb496e",
   611 => x"58a6c487",
   612 => x"ffcf4970",
   613 => x"99f8ffff",
   614 => x"87d602a9",
   615 => x"89c24970",
   616 => x"bfc0e0c2",
   617 => x"e0e4c291",
   618 => x"807148bf",
   619 => x"fc58a6c8",
   620 => x"48c087e1",
   621 => x"d0f08ef4",
   622 => x"1e731e87",
   623 => x"496a4a71",
   624 => x"7a7181c1",
   625 => x"bfc4e0c2",
   626 => x"87cb0599",
   627 => x"6b4ba2c8",
   628 => x"87fdf949",
   629 => x"c17b4970",
   630 => x"87f1ef48",
   631 => x"711e731e",
   632 => x"e0e4c24b",
   633 => x"a3c849bf",
   634 => x"c24a6a4a",
   635 => x"c0e0c28a",
   636 => x"a17292bf",
   637 => x"c4e0c249",
   638 => x"9a6b4abf",
   639 => x"c849a172",
   640 => x"e8711e66",
   641 => x"86c487fd",
   642 => x"c4059870",
   643 => x"c248c087",
   644 => x"ee48c187",
   645 => x"5e0e87f7",
   646 => x"710e5c5b",
   647 => x"724bc04a",
   648 => x"e0c0029a",
   649 => x"49a2da87",
   650 => x"c24b699f",
   651 => x"02bfc8e0",
   652 => x"a2d487cf",
   653 => x"49699f49",
   654 => x"ffffc04c",
   655 => x"c234d09c",
   656 => x"744cc087",
   657 => x"029b73b3",
   658 => x"c24a87df",
   659 => x"c0e0c28a",
   660 => x"c29249bf",
   661 => x"48bfe0e4",
   662 => x"e5c28072",
   663 => x"487158c0",
   664 => x"e0c230c4",
   665 => x"e9c058d0",
   666 => x"e4e4c287",
   667 => x"e4c24bbf",
   668 => x"e4c248fc",
   669 => x"c278bfe8",
   670 => x"02bfc8e0",
   671 => x"e0c287c9",
   672 => x"c449bfc0",
   673 => x"c287c731",
   674 => x"49bfece4",
   675 => x"e0c231c4",
   676 => x"e4c259d0",
   677 => x"f2ec5bfc",
   678 => x"5b5e0e87",
   679 => x"f40e5d5c",
   680 => x"9a4a7186",
   681 => x"c287de02",
   682 => x"c048fcd7",
   683 => x"f4d7c278",
   684 => x"fce4c248",
   685 => x"d7c278bf",
   686 => x"e4c248f8",
   687 => x"c078bff8",
   688 => x"c048eff1",
   689 => x"cce0c278",
   690 => x"d7c249bf",
   691 => x"714abffc",
   692 => x"cbc403aa",
   693 => x"cf497287",
   694 => x"e0c00599",
   695 => x"c0d8c287",
   696 => x"f4d7c21e",
   697 => x"d7c249bf",
   698 => x"a1c148f4",
   699 => x"d2e57178",
   700 => x"c086c487",
   701 => x"c248ebf1",
   702 => x"cc78c0d8",
   703 => x"ebf1c087",
   704 => x"e0c048bf",
   705 => x"eff1c080",
   706 => x"fcd7c258",
   707 => x"80c148bf",
   708 => x"58c0d8c2",
   709 => x"000c6b27",
   710 => x"bf97bf00",
   711 => x"c2029c4c",
   712 => x"e5c387ee",
   713 => x"e7c202ac",
   714 => x"ebf1c087",
   715 => x"a3cb4bbf",
   716 => x"cf4d1149",
   717 => x"d6c105ad",
   718 => x"df497487",
   719 => x"cd89c199",
   720 => x"d0e0c291",
   721 => x"4aa3c181",
   722 => x"a3c35112",
   723 => x"c551124a",
   724 => x"51124aa3",
   725 => x"124aa3c7",
   726 => x"4aa3c951",
   727 => x"a3ce5112",
   728 => x"d051124a",
   729 => x"51124aa3",
   730 => x"124aa3d2",
   731 => x"4aa3d451",
   732 => x"a3d65112",
   733 => x"d851124a",
   734 => x"51124aa3",
   735 => x"124aa3dc",
   736 => x"4aa3de51",
   737 => x"f1c05112",
   738 => x"78c148ef",
   739 => x"7587c1c1",
   740 => x"0599c849",
   741 => x"7587f3c0",
   742 => x"0599d049",
   743 => x"66dc87d0",
   744 => x"87cac002",
   745 => x"66dc4973",
   746 => x"0298700f",
   747 => x"f1c087dc",
   748 => x"c005bfef",
   749 => x"e0c287c6",
   750 => x"50c048d0",
   751 => x"48eff1c0",
   752 => x"f1c078c0",
   753 => x"c248bfeb",
   754 => x"f1c087dc",
   755 => x"78c048ef",
   756 => x"bfcce0c2",
   757 => x"fcd7c249",
   758 => x"aa714abf",
   759 => x"87f5fb04",
   760 => x"bffce4c2",
   761 => x"87c8c005",
   762 => x"bfc8e0c2",
   763 => x"87f4c102",
   764 => x"bff8d7c2",
   765 => x"87d9f149",
   766 => x"58fcd7c2",
   767 => x"e0c27e70",
   768 => x"c002bfc8",
   769 => x"496e87dd",
   770 => x"ffffffcf",
   771 => x"02a999f8",
   772 => x"c487c8c0",
   773 => x"78c048a6",
   774 => x"c487e6c0",
   775 => x"78c148a6",
   776 => x"6e87dec0",
   777 => x"f8ffcf49",
   778 => x"c002a999",
   779 => x"a6c887c8",
   780 => x"c078c048",
   781 => x"a6c887c5",
   782 => x"c478c148",
   783 => x"66c848a6",
   784 => x"0566c478",
   785 => x"6e87ddc0",
   786 => x"c289c249",
   787 => x"91bfc0e0",
   788 => x"bfe0e4c2",
   789 => x"c2807148",
   790 => x"c258f8d7",
   791 => x"c048fcd7",
   792 => x"87e1f978",
   793 => x"8ef448c0",
   794 => x"0087dee5",
   795 => x"00000000",
   796 => x"1e000000",
   797 => x"c348d4ff",
   798 => x"496878ff",
   799 => x"87c60299",
   800 => x"05a9fbc0",
   801 => x"487187ee",
   802 => x"5e0e4f26",
   803 => x"710e5c5b",
   804 => x"ff4bc04a",
   805 => x"ffc348d4",
   806 => x"99496878",
   807 => x"87c1c102",
   808 => x"02a9ecc0",
   809 => x"c087fac0",
   810 => x"c002a9fb",
   811 => x"66cc87f3",
   812 => x"cc03abb7",
   813 => x"0266d087",
   814 => x"097287c7",
   815 => x"c1097997",
   816 => x"02997182",
   817 => x"83c187c2",
   818 => x"c348d4ff",
   819 => x"496878ff",
   820 => x"87cd0299",
   821 => x"02a9ecc0",
   822 => x"fbc087c7",
   823 => x"cdff05a9",
   824 => x"0266d087",
   825 => x"97c087c3",
   826 => x"a9fbc07a",
   827 => x"7387c705",
   828 => x"8c0cc04c",
   829 => x"4c7387c2",
   830 => x"87c24874",
   831 => x"4c264d26",
   832 => x"4f264b26",
   833 => x"48d4ff1e",
   834 => x"6878ffc3",
   835 => x"b7f0c049",
   836 => x"87ca04a9",
   837 => x"a9b7f9c0",
   838 => x"c087c301",
   839 => x"c1c189f0",
   840 => x"ca04a9b7",
   841 => x"b7c6c187",
   842 => x"87c301a9",
   843 => x"7189f7c0",
   844 => x"0e4f2648",
   845 => x"5d5c5b5e",
   846 => x"7186f40e",
   847 => x"4bd4ff4c",
   848 => x"c37e4dc0",
   849 => x"d0ff7bff",
   850 => x"c0c848bf",
   851 => x"a6c898c0",
   852 => x"02987058",
   853 => x"d0ff87d0",
   854 => x"c0c848bf",
   855 => x"a6c898c0",
   856 => x"05987058",
   857 => x"d0ff87f0",
   858 => x"78e1c048",
   859 => x"c2fc7bd4",
   860 => x"99497087",
   861 => x"87c7c102",
   862 => x"c87bffc3",
   863 => x"786b48a6",
   864 => x"c04866c8",
   865 => x"c802a8fb",
   866 => x"d8e5c287",
   867 => x"eec002bf",
   868 => x"714dc187",
   869 => x"e6c00299",
   870 => x"a9fbc087",
   871 => x"fb87c302",
   872 => x"ffc387d1",
   873 => x"c1496b7b",
   874 => x"cc05a9c6",
   875 => x"7bffc387",
   876 => x"48a6c87b",
   877 => x"49c0786b",
   878 => x"0599714d",
   879 => x"7587daff",
   880 => x"dec1059d",
   881 => x"7bffc387",
   882 => x"ffc34a6b",
   883 => x"48a6c47b",
   884 => x"486e786b",
   885 => x"a6c480c1",
   886 => x"49a4c858",
   887 => x"c8496997",
   888 => x"da05a966",
   889 => x"49a4c987",
   890 => x"aa496997",
   891 => x"ca87d005",
   892 => x"699749a4",
   893 => x"a966c449",
   894 => x"c187c405",
   895 => x"c887d64d",
   896 => x"ecc04866",
   897 => x"87c902a8",
   898 => x"c04866c8",
   899 => x"c405a8fb",
   900 => x"c17ec087",
   901 => x"7bffc34d",
   902 => x"6b48a6c8",
   903 => x"029d7578",
   904 => x"ff87e2fe",
   905 => x"c848bfd0",
   906 => x"c898c0c0",
   907 => x"987058a6",
   908 => x"ff87d002",
   909 => x"c848bfd0",
   910 => x"c898c0c0",
   911 => x"987058a6",
   912 => x"ff87f005",
   913 => x"e0c048d0",
   914 => x"f4486e78",
   915 => x"87ecfa8e",
   916 => x"5c5b5e0e",
   917 => x"86f40e5d",
   918 => x"ff59a6c4",
   919 => x"c0c84cd0",
   920 => x"1e6e4bc0",
   921 => x"49dce5c2",
   922 => x"c487cfe9",
   923 => x"02987086",
   924 => x"c287f7c5",
   925 => x"4dbfe0e5",
   926 => x"f6fa496e",
   927 => x"58a6c887",
   928 => x"9873486c",
   929 => x"7058a6cc",
   930 => x"87cc0298",
   931 => x"9873486c",
   932 => x"7058a6c4",
   933 => x"87f40598",
   934 => x"d4ff7cc5",
   935 => x"78d5c148",
   936 => x"bfd8e5c2",
   937 => x"c481c149",
   938 => x"8ac14a66",
   939 => x"487232c6",
   940 => x"d4ffb071",
   941 => x"486c7808",
   942 => x"a6c49873",
   943 => x"02987058",
   944 => x"486c87cc",
   945 => x"a6c49873",
   946 => x"05987058",
   947 => x"7cc487f4",
   948 => x"c348d4ff",
   949 => x"486c78ff",
   950 => x"a6c49873",
   951 => x"02987058",
   952 => x"486c87cc",
   953 => x"a6c49873",
   954 => x"05987058",
   955 => x"7cc587f4",
   956 => x"c148d4ff",
   957 => x"78c178d3",
   958 => x"9873486c",
   959 => x"7058a6c4",
   960 => x"87cc0298",
   961 => x"9873486c",
   962 => x"7058a6c4",
   963 => x"87f40598",
   964 => x"9d757cc4",
   965 => x"87d0c202",
   966 => x"7ec0d8c2",
   967 => x"dce5c21e",
   968 => x"87f8ea49",
   969 => x"987086c4",
   970 => x"c087c505",
   971 => x"87fcc248",
   972 => x"adb7c0c8",
   973 => x"4a87c404",
   974 => x"7587c48d",
   975 => x"6c4dc04a",
   976 => x"c8987348",
   977 => x"987058a6",
   978 => x"6c87cc02",
   979 => x"c8987348",
   980 => x"987058a6",
   981 => x"cd87f405",
   982 => x"48d4ff7c",
   983 => x"7278d4c1",
   984 => x"718ac149",
   985 => x"87d90299",
   986 => x"48bf976e",
   987 => x"7808d4ff",
   988 => x"80c1486e",
   989 => x"7258a6c4",
   990 => x"718ac149",
   991 => x"e7ff0599",
   992 => x"73486c87",
   993 => x"58a6c498",
   994 => x"cc029870",
   995 => x"73486c87",
   996 => x"58a6c498",
   997 => x"f4059870",
   998 => x"c27cc487",
   999 => x"e849dce5",
  1000 => x"9d7587d7",
  1001 => x"87f0fd05",
  1002 => x"9873486c",
  1003 => x"7058a6c4",
  1004 => x"87cd0298",
  1005 => x"9873486c",
  1006 => x"7058a6c4",
  1007 => x"f3ff0598",
  1008 => x"ff7cc587",
  1009 => x"d3c148d4",
  1010 => x"6c78c078",
  1011 => x"c4987348",
  1012 => x"987058a6",
  1013 => x"6c87cd02",
  1014 => x"c4987348",
  1015 => x"987058a6",
  1016 => x"87f3ff05",
  1017 => x"48c17cc4",
  1018 => x"48c087c2",
  1019 => x"cbf48ef4",
  1020 => x"5b5e0e87",
  1021 => x"1e0e5d5c",
  1022 => x"4cc04b71",
  1023 => x"04abb74d",
  1024 => x"c087e9c0",
  1025 => x"751ef3f4",
  1026 => x"87c4029d",
  1027 => x"87c24ac0",
  1028 => x"49724ac1",
  1029 => x"c487c2ea",
  1030 => x"c158a686",
  1031 => x"c2056e84",
  1032 => x"c14c7387",
  1033 => x"acb77385",
  1034 => x"87d7ff06",
  1035 => x"f326486e",
  1036 => x"5e0e87ca",
  1037 => x"0e5d5c5b",
  1038 => x"494c711e",
  1039 => x"bfece5c2",
  1040 => x"87edfe81",
  1041 => x"029d4d70",
  1042 => x"c287fcc0",
  1043 => x"754bd0e0",
  1044 => x"ff49cb4a",
  1045 => x"7487c9c1",
  1046 => x"c291de49",
  1047 => x"7148c0e6",
  1048 => x"58a6c480",
  1049 => x"48d7c2c1",
  1050 => x"a1c8496e",
  1051 => x"7141204a",
  1052 => x"87f905aa",
  1053 => x"51105110",
  1054 => x"49745110",
  1055 => x"87eec5c1",
  1056 => x"49d0e0c2",
  1057 => x"c187c9f7",
  1058 => x"c149d0e4",
  1059 => x"c187f6c7",
  1060 => x"2687d2c8",
  1061 => x"4c87e5f1",
  1062 => x"6964616f",
  1063 => x"2e2e676e",
  1064 => x"2080002e",
  1065 => x"6b636142",
  1066 => x"616f4c00",
  1067 => x"2e2a2064",
  1068 => x"203a0020",
  1069 => x"42208000",
  1070 => x"006b6361",
  1071 => x"78452080",
  1072 => x"53007469",
  1073 => x"6e492044",
  1074 => x"2e2e7469",
  1075 => x"004b4f00",
  1076 => x"544f4f42",
  1077 => x"20202020",
  1078 => x"004d4f52",
  1079 => x"711e731e",
  1080 => x"e5c2494b",
  1081 => x"fc81bfec",
  1082 => x"4a7087c7",
  1083 => x"87c4029a",
  1084 => x"87e2e449",
  1085 => x"48ece5c2",
  1086 => x"497378c0",
  1087 => x"ef87e9c1",
  1088 => x"731e87fe",
  1089 => x"c44b711e",
  1090 => x"c1024aa3",
  1091 => x"8ac187c8",
  1092 => x"8a87dc02",
  1093 => x"87f1c002",
  1094 => x"c4c1058a",
  1095 => x"ece5c287",
  1096 => x"fcc002bf",
  1097 => x"88c14887",
  1098 => x"58f0e5c2",
  1099 => x"c287f2c0",
  1100 => x"49bfece5",
  1101 => x"e5c289d0",
  1102 => x"b7c059f0",
  1103 => x"e0c003a9",
  1104 => x"ece5c287",
  1105 => x"d878c048",
  1106 => x"ece5c287",
  1107 => x"80c148bf",
  1108 => x"58f0e5c2",
  1109 => x"e5c287cb",
  1110 => x"d048bfec",
  1111 => x"f0e5c280",
  1112 => x"c3497358",
  1113 => x"87d8ee87",
  1114 => x"5c5b5e0e",
  1115 => x"86f00e5d",
  1116 => x"c259a6d0",
  1117 => x"c04dc0d8",
  1118 => x"48a6c44c",
  1119 => x"e5c278c0",
  1120 => x"c048bfec",
  1121 => x"c106a8b7",
  1122 => x"d8c287c1",
  1123 => x"029848c0",
  1124 => x"c087f8c0",
  1125 => x"c81ef3f4",
  1126 => x"87c70266",
  1127 => x"c048a6c4",
  1128 => x"c487c578",
  1129 => x"78c148a6",
  1130 => x"e34966c4",
  1131 => x"86c487eb",
  1132 => x"84c14d70",
  1133 => x"c14866c4",
  1134 => x"58a6c880",
  1135 => x"bfece5c2",
  1136 => x"c603acb7",
  1137 => x"059d7587",
  1138 => x"c087c8ff",
  1139 => x"029d754c",
  1140 => x"c087e3c3",
  1141 => x"c81ef3f4",
  1142 => x"87c70266",
  1143 => x"c048a6cc",
  1144 => x"cc87c578",
  1145 => x"78c148a6",
  1146 => x"e24966cc",
  1147 => x"86c487eb",
  1148 => x"026e58a6",
  1149 => x"4987ebc2",
  1150 => x"699781cb",
  1151 => x"0299d049",
  1152 => x"c187d9c1",
  1153 => x"744bdcc3",
  1154 => x"c191cc49",
  1155 => x"c881d0e4",
  1156 => x"7a734aa1",
  1157 => x"ffc381c1",
  1158 => x"de497451",
  1159 => x"c0e6c291",
  1160 => x"c285714d",
  1161 => x"c17d97c1",
  1162 => x"e0c049a5",
  1163 => x"d0e0c251",
  1164 => x"d202bf97",
  1165 => x"c284c187",
  1166 => x"e0c24ba5",
  1167 => x"49db4ad0",
  1168 => x"87dcf9fe",
  1169 => x"cd87dbc1",
  1170 => x"51c049a5",
  1171 => x"a5c284c1",
  1172 => x"cb4a6e4b",
  1173 => x"c7f9fe49",
  1174 => x"87c6c187",
  1175 => x"91cc4974",
  1176 => x"81d0e4c1",
  1177 => x"c0c181c8",
  1178 => x"e0c279f2",
  1179 => x"02bf97d0",
  1180 => x"497487d8",
  1181 => x"84c191de",
  1182 => x"4bc0e6c2",
  1183 => x"e0c28371",
  1184 => x"49dd4ad0",
  1185 => x"87d8f8fe",
  1186 => x"4b7487d8",
  1187 => x"e6c293de",
  1188 => x"a3cb83c0",
  1189 => x"c151c049",
  1190 => x"4a6e7384",
  1191 => x"f7fe49cb",
  1192 => x"66c487fe",
  1193 => x"c880c148",
  1194 => x"b7c758a6",
  1195 => x"c5c003ac",
  1196 => x"fc056e87",
  1197 => x"b7c787dd",
  1198 => x"d3c003ac",
  1199 => x"de497487",
  1200 => x"c0e6c291",
  1201 => x"c151c081",
  1202 => x"acb7c784",
  1203 => x"87edff04",
  1204 => x"48e5e5c1",
  1205 => x"e5c150c0",
  1206 => x"50c248e4",
  1207 => x"48ece5c1",
  1208 => x"78ceccc1",
  1209 => x"48e8e5c1",
  1210 => x"78e2c2c1",
  1211 => x"48f8e5c1",
  1212 => x"78c2c4c1",
  1213 => x"c04966cc",
  1214 => x"f087f3fb",
  1215 => x"87fce78e",
  1216 => x"c24a711e",
  1217 => x"725adce5",
  1218 => x"87dcf949",
  1219 => x"711e4f26",
  1220 => x"91cc494a",
  1221 => x"81d0e4c1",
  1222 => x"481181c1",
  1223 => x"58d8e5c2",
  1224 => x"49a2f0c0",
  1225 => x"87c8f6fe",
  1226 => x"ddd549c0",
  1227 => x"0e4f2687",
  1228 => x"5d5c5b5e",
  1229 => x"7186f00e",
  1230 => x"91cc494c",
  1231 => x"81d0e4c1",
  1232 => x"c47ea1c3",
  1233 => x"e5c248a6",
  1234 => x"6e78bfd0",
  1235 => x"c44abf97",
  1236 => x"2b724b66",
  1237 => x"124aa1c1",
  1238 => x"58a6cc48",
  1239 => x"83c19b70",
  1240 => x"699781c2",
  1241 => x"04abb749",
  1242 => x"4bc087c2",
  1243 => x"4abf976e",
  1244 => x"724966c8",
  1245 => x"c4b9ff31",
  1246 => x"4d739966",
  1247 => x"b5713572",
  1248 => x"5dd4e5c2",
  1249 => x"c348d4ff",
  1250 => x"d0ff78ff",
  1251 => x"c0c848bf",
  1252 => x"a6d098c0",
  1253 => x"02987058",
  1254 => x"d0ff87d0",
  1255 => x"c0c848bf",
  1256 => x"a6c498c0",
  1257 => x"05987058",
  1258 => x"d0ff87f0",
  1259 => x"78e1c048",
  1260 => x"de48d4ff",
  1261 => x"7d0d7078",
  1262 => x"c848750d",
  1263 => x"d4ff28b7",
  1264 => x"48757808",
  1265 => x"ff28b7d0",
  1266 => x"757808d4",
  1267 => x"28b7d848",
  1268 => x"7808d4ff",
  1269 => x"48bfd0ff",
  1270 => x"98c0c0c8",
  1271 => x"7058a6c4",
  1272 => x"87d00298",
  1273 => x"48bfd0ff",
  1274 => x"98c0c0c8",
  1275 => x"7058a6c4",
  1276 => x"87f00598",
  1277 => x"c048d0ff",
  1278 => x"1ec778e0",
  1279 => x"e4c11ec0",
  1280 => x"e5c21ed0",
  1281 => x"c149bfd4",
  1282 => x"497487e1",
  1283 => x"87def7c0",
  1284 => x"e7e38ee4",
  1285 => x"1e731e87",
  1286 => x"fc494b71",
  1287 => x"497387d1",
  1288 => x"e387ccfc",
  1289 => x"731e87da",
  1290 => x"c24b711e",
  1291 => x"d5024aa3",
  1292 => x"058ac187",
  1293 => x"e5c287db",
  1294 => x"d402bfe8",
  1295 => x"88c14887",
  1296 => x"58ece5c2",
  1297 => x"e5c287cb",
  1298 => x"c148bfe8",
  1299 => x"ece5c280",
  1300 => x"c01ec758",
  1301 => x"d0e4c11e",
  1302 => x"d4e5c21e",
  1303 => x"87cb49bf",
  1304 => x"f6c04973",
  1305 => x"8ef487c8",
  1306 => x"0e87d5e2",
  1307 => x"5d5c5b5e",
  1308 => x"86d8ff0e",
  1309 => x"c859a6dc",
  1310 => x"78c048a6",
  1311 => x"78c080c4",
  1312 => x"c280c44d",
  1313 => x"78bfe8e5",
  1314 => x"c348d4ff",
  1315 => x"d0ff78ff",
  1316 => x"c0c848bf",
  1317 => x"a6c498c0",
  1318 => x"02987058",
  1319 => x"d0ff87d0",
  1320 => x"c0c848bf",
  1321 => x"a6c498c0",
  1322 => x"05987058",
  1323 => x"d0ff87f0",
  1324 => x"78e1c048",
  1325 => x"d448d4ff",
  1326 => x"f6deff78",
  1327 => x"48d4ff87",
  1328 => x"d478ffc3",
  1329 => x"d4ff48a6",
  1330 => x"66d478bf",
  1331 => x"a8fbc048",
  1332 => x"87d3c102",
  1333 => x"4a66f8c0",
  1334 => x"7e6a82c4",
  1335 => x"c2c11e72",
  1336 => x"66c448e9",
  1337 => x"4aa1c849",
  1338 => x"aa714120",
  1339 => x"1087f905",
  1340 => x"c04a2651",
  1341 => x"c84966f8",
  1342 => x"c0ccc181",
  1343 => x"c7496a79",
  1344 => x"5166d481",
  1345 => x"1ed81ec1",
  1346 => x"81c8496a",
  1347 => x"87faddff",
  1348 => x"66d086c8",
  1349 => x"a8b7c048",
  1350 => x"c187c401",
  1351 => x"d087c84d",
  1352 => x"88c14866",
  1353 => x"d458a6d4",
  1354 => x"f4ca0266",
  1355 => x"66c0c187",
  1356 => x"ca03adb7",
  1357 => x"d4ff87eb",
  1358 => x"78ffc348",
  1359 => x"ff48a6d4",
  1360 => x"d478bfd4",
  1361 => x"c6c14866",
  1362 => x"58a6c488",
  1363 => x"c0029870",
  1364 => x"c94887e6",
  1365 => x"58a6c488",
  1366 => x"c4029870",
  1367 => x"c14887d5",
  1368 => x"58a6c488",
  1369 => x"c1029870",
  1370 => x"c44887e3",
  1371 => x"7058a688",
  1372 => x"fec30298",
  1373 => x"87d3c987",
  1374 => x"c10566d8",
  1375 => x"d4ff87c5",
  1376 => x"78ffc348",
  1377 => x"1eca1ec0",
  1378 => x"93cc4b75",
  1379 => x"8366c0c1",
  1380 => x"6c4ca3c4",
  1381 => x"f1dbff49",
  1382 => x"de1ec187",
  1383 => x"ff496c1e",
  1384 => x"d087e7db",
  1385 => x"49a3c886",
  1386 => x"79c0ccc1",
  1387 => x"adb766d0",
  1388 => x"c187c504",
  1389 => x"87dac885",
  1390 => x"c14866d0",
  1391 => x"58a6d488",
  1392 => x"ff87cfc8",
  1393 => x"d887ecda",
  1394 => x"c5c858a6",
  1395 => x"f3dcff87",
  1396 => x"58a6cc87",
  1397 => x"a8b766cc",
  1398 => x"cc87c606",
  1399 => x"66c848a6",
  1400 => x"dfdcff78",
  1401 => x"a8ecc087",
  1402 => x"87c7c205",
  1403 => x"c10566d8",
  1404 => x"497587f7",
  1405 => x"f8c091cc",
  1406 => x"a1c48166",
  1407 => x"c14c6a4a",
  1408 => x"66c84aa1",
  1409 => x"7997c252",
  1410 => x"ccc181c8",
  1411 => x"d4ff79ce",
  1412 => x"78ffc348",
  1413 => x"ff48a6d4",
  1414 => x"d478bfd4",
  1415 => x"e8c00266",
  1416 => x"fbc04887",
  1417 => x"e0c002a8",
  1418 => x"9766d487",
  1419 => x"ff84c17c",
  1420 => x"ffc348d4",
  1421 => x"48a6d478",
  1422 => x"78bfd4ff",
  1423 => x"c80266d4",
  1424 => x"fbc04887",
  1425 => x"e0ff05a8",
  1426 => x"54e0c087",
  1427 => x"c054c1c2",
  1428 => x"66d07c97",
  1429 => x"c504adb7",
  1430 => x"c585c187",
  1431 => x"66d087f4",
  1432 => x"d488c148",
  1433 => x"e9c558a6",
  1434 => x"c6d8ff87",
  1435 => x"58a6d887",
  1436 => x"c887dfc5",
  1437 => x"66d84866",
  1438 => x"c4c505a8",
  1439 => x"48a6dc87",
  1440 => x"d9ff78c0",
  1441 => x"a6d887fe",
  1442 => x"f7d9ff58",
  1443 => x"a6e4c087",
  1444 => x"a8ecc058",
  1445 => x"87cac005",
  1446 => x"48a6e0c0",
  1447 => x"c07866d4",
  1448 => x"d4ff87c6",
  1449 => x"78ffc348",
  1450 => x"91cc4975",
  1451 => x"4866f8c0",
  1452 => x"a6c48071",
  1453 => x"c3496e58",
  1454 => x"5166d481",
  1455 => x"4966e0c0",
  1456 => x"66d481c1",
  1457 => x"7148c189",
  1458 => x"c1497030",
  1459 => x"c14a6e89",
  1460 => x"97097282",
  1461 => x"486e0979",
  1462 => x"e5c250c2",
  1463 => x"d449bfd0",
  1464 => x"9729b766",
  1465 => x"71484a6a",
  1466 => x"a6e8c098",
  1467 => x"c4486e58",
  1468 => x"58a6c880",
  1469 => x"4cbf66c4",
  1470 => x"c84866d8",
  1471 => x"c002a866",
  1472 => x"e0c087c9",
  1473 => x"78c048a6",
  1474 => x"c087c6c0",
  1475 => x"c148a6e0",
  1476 => x"66e0c078",
  1477 => x"1ee0c01e",
  1478 => x"d5ff4974",
  1479 => x"86c887ec",
  1480 => x"c058a6d8",
  1481 => x"c106a8b7",
  1482 => x"66d487da",
  1483 => x"bf66c484",
  1484 => x"81e0c049",
  1485 => x"c14b8974",
  1486 => x"714af2c2",
  1487 => x"87e0e5fe",
  1488 => x"66dc84c2",
  1489 => x"c080c148",
  1490 => x"c058a6e0",
  1491 => x"c14966e4",
  1492 => x"02a97081",
  1493 => x"c087c9c0",
  1494 => x"c048a6e0",
  1495 => x"87c6c078",
  1496 => x"48a6e0c0",
  1497 => x"e0c078c1",
  1498 => x"66c81e66",
  1499 => x"e0c049bf",
  1500 => x"71897481",
  1501 => x"ff49741e",
  1502 => x"c887cfd4",
  1503 => x"a8b7c086",
  1504 => x"87fefe01",
  1505 => x"c00266dc",
  1506 => x"496e87d2",
  1507 => x"66dc81c2",
  1508 => x"c8496e51",
  1509 => x"efccc181",
  1510 => x"87cdc079",
  1511 => x"81c2496e",
  1512 => x"c8496e51",
  1513 => x"d5d0c181",
  1514 => x"b766d079",
  1515 => x"c5c004ad",
  1516 => x"c085c187",
  1517 => x"66d087dc",
  1518 => x"d488c148",
  1519 => x"d1c058a6",
  1520 => x"eed2ff87",
  1521 => x"58a6d887",
  1522 => x"ff87c7c0",
  1523 => x"d887e4d2",
  1524 => x"66d458a6",
  1525 => x"87c9c002",
  1526 => x"b766c0c1",
  1527 => x"d5f504ad",
  1528 => x"adb7c787",
  1529 => x"87dcc003",
  1530 => x"91cc4975",
  1531 => x"8166f8c0",
  1532 => x"6a4aa1c4",
  1533 => x"c852c04a",
  1534 => x"c179c081",
  1535 => x"adb7c785",
  1536 => x"87e4ff04",
  1537 => x"c00266d8",
  1538 => x"f8c087eb",
  1539 => x"d4c14966",
  1540 => x"66f8c081",
  1541 => x"82d5c14a",
  1542 => x"51c252c0",
  1543 => x"4966f8c0",
  1544 => x"c181dcc1",
  1545 => x"c079cecc",
  1546 => x"c14966f8",
  1547 => x"c2c181d8",
  1548 => x"d6c079f5",
  1549 => x"66f8c087",
  1550 => x"81d8c149",
  1551 => x"79fcc2c1",
  1552 => x"4966f8c0",
  1553 => x"c281dcc1",
  1554 => x"c179e5ca",
  1555 => x"c04ae6d0",
  1556 => x"c14966f8",
  1557 => x"797281e8",
  1558 => x"48bfd0ff",
  1559 => x"98c0c0c8",
  1560 => x"7058a6c4",
  1561 => x"d1c00298",
  1562 => x"bfd0ff87",
  1563 => x"c0c0c848",
  1564 => x"58a6c498",
  1565 => x"ff059870",
  1566 => x"d0ff87ef",
  1567 => x"78e0c048",
  1568 => x"ff4866cc",
  1569 => x"d1ff8ed8",
  1570 => x"c71e87f2",
  1571 => x"c11ec01e",
  1572 => x"c21ed0e4",
  1573 => x"49bfd4e5",
  1574 => x"c187d0ef",
  1575 => x"c049d0e4",
  1576 => x"f487e2e7",
  1577 => x"1e4f268e",
  1578 => x"c287c6ca",
  1579 => x"c048f0e5",
  1580 => x"48d4ff50",
  1581 => x"c178ffc3",
  1582 => x"fe49c3c3",
  1583 => x"fe87fdde",
  1584 => x"7087c8e8",
  1585 => x"87cd0298",
  1586 => x"87c5f4fe",
  1587 => x"c4029870",
  1588 => x"c24ac187",
  1589 => x"724ac087",
  1590 => x"87c8029a",
  1591 => x"49cdc3c1",
  1592 => x"87d8defe",
  1593 => x"bfc0d7c2",
  1594 => x"e3d5ff49",
  1595 => x"e8e5c287",
  1596 => x"c278c048",
  1597 => x"c048d4e5",
  1598 => x"cdfe4978",
  1599 => x"87ddc387",
  1600 => x"c087c2c9",
  1601 => x"ff87ede6",
  1602 => x"4f2687f6",
  1603 => x"000010d0",
  1604 => x"00000002",
  1605 => x"00002980",
  1606 => x"00001032",
  1607 => x"00000002",
  1608 => x"0000299e",
  1609 => x"00001032",
  1610 => x"00000002",
  1611 => x"000029bc",
  1612 => x"00001032",
  1613 => x"00000002",
  1614 => x"000029da",
  1615 => x"00001032",
  1616 => x"00000002",
  1617 => x"000029f8",
  1618 => x"00001032",
  1619 => x"00000002",
  1620 => x"00002a16",
  1621 => x"00001032",
  1622 => x"00000002",
  1623 => x"00002a34",
  1624 => x"00001032",
  1625 => x"00000002",
  1626 => x"00000000",
  1627 => x"0000130e",
  1628 => x"00000000",
  1629 => x"00000000",
  1630 => x"00001102",
  1631 => x"d5c11e1e",
  1632 => x"58a6c487",
  1633 => x"1e4f2626",
  1634 => x"f0fe4a71",
  1635 => x"cd78c048",
  1636 => x"c10a7a0a",
  1637 => x"fe49dde6",
  1638 => x"2687e1db",
  1639 => x"7465534f",
  1640 => x"6e616820",
  1641 => x"72656c64",
  1642 => x"6e49000a",
  1643 => x"746e6920",
  1644 => x"75727265",
  1645 => x"63207470",
  1646 => x"74736e6f",
  1647 => x"74637572",
  1648 => x"000a726f",
  1649 => x"eae6c11e",
  1650 => x"efdafe49",
  1651 => x"fce5c187",
  1652 => x"87f3fe49",
  1653 => x"fe1e4f26",
  1654 => x"2648bff0",
  1655 => x"f0fe1e4f",
  1656 => x"2678c148",
  1657 => x"f0fe1e4f",
  1658 => x"2678c048",
  1659 => x"4a711e4f",
  1660 => x"a2c47ac0",
  1661 => x"c879c049",
  1662 => x"79c049a2",
  1663 => x"c049a2cc",
  1664 => x"0e4f2679",
  1665 => x"0e5c5b5e",
  1666 => x"4c7186f8",
  1667 => x"cc49a4c8",
  1668 => x"486b4ba4",
  1669 => x"a6c480c1",
  1670 => x"c898cf58",
  1671 => x"486958a6",
  1672 => x"05a866c4",
  1673 => x"486b87d4",
  1674 => x"a6c480c1",
  1675 => x"c898cf58",
  1676 => x"486958a6",
  1677 => x"02a866c4",
  1678 => x"e8fe87ec",
  1679 => x"a4d0c187",
  1680 => x"c4486b49",
  1681 => x"58a6c490",
  1682 => x"66d48170",
  1683 => x"c1486b79",
  1684 => x"58a6c880",
  1685 => x"7b7098cf",
  1686 => x"fd87d2c1",
  1687 => x"8ef887ff",
  1688 => x"4d2687c2",
  1689 => x"4b264c26",
  1690 => x"5e0e4f26",
  1691 => x"0e5d5c5b",
  1692 => x"4d7186f8",
  1693 => x"6d4ca5c4",
  1694 => x"05a86c48",
  1695 => x"48ff87c5",
  1696 => x"fd87e5c0",
  1697 => x"a5d087df",
  1698 => x"c4486c4b",
  1699 => x"58a6c490",
  1700 => x"4b6b8370",
  1701 => x"6c9bffc3",
  1702 => x"c880c148",
  1703 => x"98cf58a6",
  1704 => x"f8fc7c70",
  1705 => x"48497387",
  1706 => x"f5fe8ef8",
  1707 => x"1e731e87",
  1708 => x"f0fc86f8",
  1709 => x"4bbfe087",
  1710 => x"c0e0c049",
  1711 => x"e7c00299",
  1712 => x"c34a7387",
  1713 => x"e9c29aff",
  1714 => x"c448bfd2",
  1715 => x"58a6c490",
  1716 => x"49e2e9c2",
  1717 => x"79728170",
  1718 => x"bfd2e9c2",
  1719 => x"c880c148",
  1720 => x"98cf58a6",
  1721 => x"58d6e9c2",
  1722 => x"c0d04973",
  1723 => x"f2c00299",
  1724 => x"dae9c287",
  1725 => x"e9c248bf",
  1726 => x"02a8bfde",
  1727 => x"c287e4c0",
  1728 => x"48bfdae9",
  1729 => x"a6c490c4",
  1730 => x"e2eac258",
  1731 => x"e0817049",
  1732 => x"c2786948",
  1733 => x"48bfdae9",
  1734 => x"a6c880c1",
  1735 => x"c298cf58",
  1736 => x"fa58dee9",
  1737 => x"a6c487f0",
  1738 => x"87f1fa58",
  1739 => x"f5fc8ef8",
  1740 => x"e9c21e87",
  1741 => x"f4fa49d2",
  1742 => x"edeac187",
  1743 => x"87c7f949",
  1744 => x"2687f5c3",
  1745 => x"1e731e4f",
  1746 => x"49d2e9c2",
  1747 => x"7087dbfc",
  1748 => x"aab7c04a",
  1749 => x"87ccc204",
  1750 => x"05aaf0c3",
  1751 => x"efc187c9",
  1752 => x"78c148f0",
  1753 => x"c387edc1",
  1754 => x"c905aae0",
  1755 => x"f4efc187",
  1756 => x"c178c148",
  1757 => x"efc187de",
  1758 => x"c602bff4",
  1759 => x"a2c0c287",
  1760 => x"7287c24b",
  1761 => x"f0efc14b",
  1762 => x"e0c002bf",
  1763 => x"c4497387",
  1764 => x"c19129b7",
  1765 => x"7381f8ef",
  1766 => x"c29acf4a",
  1767 => x"7248c192",
  1768 => x"ff4a7030",
  1769 => x"694872ba",
  1770 => x"db797098",
  1771 => x"c4497387",
  1772 => x"c19129b7",
  1773 => x"7381f8ef",
  1774 => x"c29acf4a",
  1775 => x"7248c392",
  1776 => x"484a7030",
  1777 => x"7970b069",
  1778 => x"48f4efc1",
  1779 => x"efc178c0",
  1780 => x"78c048f0",
  1781 => x"49d2e9c2",
  1782 => x"7087cffa",
  1783 => x"aab7c04a",
  1784 => x"87f4fd03",
  1785 => x"87c448c0",
  1786 => x"4c264d26",
  1787 => x"4f264b26",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"724ac01e",
  1807 => x"c191c449",
  1808 => x"c081f8ef",
  1809 => x"d082c179",
  1810 => x"ee04aab7",
  1811 => x"0e4f2687",
  1812 => x"5d5c5b5e",
  1813 => x"f64d710e",
  1814 => x"4a7587cb",
  1815 => x"922ab7c4",
  1816 => x"82f8efc1",
  1817 => x"9ccf4c75",
  1818 => x"496a94c2",
  1819 => x"c32b744b",
  1820 => x"7448c29b",
  1821 => x"ff4c7030",
  1822 => x"714874bc",
  1823 => x"f57a7098",
  1824 => x"487387db",
  1825 => x"1e87e1fd",
  1826 => x"bfd0ff1e",
  1827 => x"c0c0c848",
  1828 => x"58a6c498",
  1829 => x"d0029870",
  1830 => x"bfd0ff87",
  1831 => x"c0c0c848",
  1832 => x"58a6c498",
  1833 => x"f0059870",
  1834 => x"48d0ff87",
  1835 => x"7178e1c4",
  1836 => x"08d4ff48",
  1837 => x"4866c878",
  1838 => x"7808d4ff",
  1839 => x"1e4f2626",
  1840 => x"c84a711e",
  1841 => x"721e4966",
  1842 => x"87fbfe49",
  1843 => x"d0ff86c4",
  1844 => x"c0c848bf",
  1845 => x"a6c498c0",
  1846 => x"02987058",
  1847 => x"d0ff87d0",
  1848 => x"c0c848bf",
  1849 => x"a6c498c0",
  1850 => x"05987058",
  1851 => x"d0ff87f0",
  1852 => x"78e0c048",
  1853 => x"1e4f2626",
  1854 => x"4b711e73",
  1855 => x"731e66c8",
  1856 => x"a2e0c14a",
  1857 => x"87f7fe49",
  1858 => x"2687c426",
  1859 => x"264c264d",
  1860 => x"1e4f264b",
  1861 => x"bfd0ff1e",
  1862 => x"c0c0c848",
  1863 => x"58a6c498",
  1864 => x"d0029870",
  1865 => x"bfd0ff87",
  1866 => x"c0c0c848",
  1867 => x"58a6c498",
  1868 => x"f0059870",
  1869 => x"48d0ff87",
  1870 => x"7178c9c4",
  1871 => x"08d4ff48",
  1872 => x"4f262678",
  1873 => x"4a711e1e",
  1874 => x"87c7ff49",
  1875 => x"48bfd0ff",
  1876 => x"98c0c0c8",
  1877 => x"7058a6c4",
  1878 => x"87d00298",
  1879 => x"48bfd0ff",
  1880 => x"98c0c0c8",
  1881 => x"7058a6c4",
  1882 => x"87f00598",
  1883 => x"c848d0ff",
  1884 => x"4f262678",
  1885 => x"1e1e731e",
  1886 => x"ebc24b71",
  1887 => x"c302bfee",
  1888 => x"87ccc387",
  1889 => x"48bfd0ff",
  1890 => x"98c0c0c8",
  1891 => x"7058a6c4",
  1892 => x"87d00298",
  1893 => x"48bfd0ff",
  1894 => x"98c0c0c8",
  1895 => x"7058a6c4",
  1896 => x"87f00598",
  1897 => x"c448d0ff",
  1898 => x"487378c9",
  1899 => x"ffb0e0c0",
  1900 => x"c27808d4",
  1901 => x"c048e2eb",
  1902 => x"0266cc78",
  1903 => x"ffc387c5",
  1904 => x"c087c249",
  1905 => x"eaebc249",
  1906 => x"0266d059",
  1907 => x"d5c587c6",
  1908 => x"87c44ad5",
  1909 => x"4affffcf",
  1910 => x"5aeeebc2",
  1911 => x"48eeebc2",
  1912 => x"c42678c1",
  1913 => x"264d2687",
  1914 => x"264b264c",
  1915 => x"5b5e0e4f",
  1916 => x"710e5d5c",
  1917 => x"eaebc24a",
  1918 => x"9a724cbf",
  1919 => x"4987cb02",
  1920 => x"f6c191c8",
  1921 => x"83714bee",
  1922 => x"fac187c4",
  1923 => x"4dc04bee",
  1924 => x"99744913",
  1925 => x"bfe6ebc2",
  1926 => x"ffb87148",
  1927 => x"c17808d4",
  1928 => x"c8852cb7",
  1929 => x"e704adb7",
  1930 => x"e2ebc287",
  1931 => x"80c848bf",
  1932 => x"58e6ebc2",
  1933 => x"1e87eefe",
  1934 => x"4b711e73",
  1935 => x"029a4a13",
  1936 => x"497287cb",
  1937 => x"1387e6fe",
  1938 => x"f5059a4a",
  1939 => x"87d9fe87",
  1940 => x"ebc21e1e",
  1941 => x"c249bfe2",
  1942 => x"c148e2eb",
  1943 => x"c0c478a1",
  1944 => x"db03a9b7",
  1945 => x"48d4ff87",
  1946 => x"bfe6ebc2",
  1947 => x"e2ebc278",
  1948 => x"ebc249bf",
  1949 => x"a1c148e2",
  1950 => x"b7c0c478",
  1951 => x"87e504a9",
  1952 => x"48bfd0ff",
  1953 => x"98c0c0c8",
  1954 => x"7058a6c4",
  1955 => x"87d00298",
  1956 => x"48bfd0ff",
  1957 => x"98c0c0c8",
  1958 => x"7058a6c4",
  1959 => x"87f00598",
  1960 => x"c848d0ff",
  1961 => x"eeebc278",
  1962 => x"2678c048",
  1963 => x"00004f26",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"005f5f00",
  1967 => x"03000000",
  1968 => x"03030003",
  1969 => x"7f140000",
  1970 => x"7f7f147f",
  1971 => x"24000014",
  1972 => x"3a6b6b2e",
  1973 => x"6a4c0012",
  1974 => x"566c1836",
  1975 => x"7e300032",
  1976 => x"3a77594f",
  1977 => x"00004068",
  1978 => x"00030704",
  1979 => x"00000000",
  1980 => x"41633e1c",
  1981 => x"00000000",
  1982 => x"1c3e6341",
  1983 => x"2a080000",
  1984 => x"3e1c1c3e",
  1985 => x"0800082a",
  1986 => x"083e3e08",
  1987 => x"00000008",
  1988 => x"0060e080",
  1989 => x"08000000",
  1990 => x"08080808",
  1991 => x"00000008",
  1992 => x"00606000",
  1993 => x"60400000",
  1994 => x"060c1830",
  1995 => x"3e000103",
  1996 => x"7f4d597f",
  1997 => x"0400003e",
  1998 => x"007f7f06",
  1999 => x"42000000",
  2000 => x"4f597163",
  2001 => x"22000046",
  2002 => x"7f494963",
  2003 => x"1c180036",
  2004 => x"7f7f1316",
  2005 => x"27000010",
  2006 => x"7d454567",
  2007 => x"3c000039",
  2008 => x"79494b7e",
  2009 => x"01000030",
  2010 => x"0f797101",
  2011 => x"36000007",
  2012 => x"7f49497f",
  2013 => x"06000036",
  2014 => x"3f69494f",
  2015 => x"0000001e",
  2016 => x"00666600",
  2017 => x"00000000",
  2018 => x"0066e680",
  2019 => x"08000000",
  2020 => x"22141408",
  2021 => x"14000022",
  2022 => x"14141414",
  2023 => x"22000014",
  2024 => x"08141422",
  2025 => x"02000008",
  2026 => x"0f595103",
  2027 => x"7f3e0006",
  2028 => x"1f555d41",
  2029 => x"7e00001e",
  2030 => x"7f09097f",
  2031 => x"7f00007e",
  2032 => x"7f49497f",
  2033 => x"1c000036",
  2034 => x"4141633e",
  2035 => x"7f000041",
  2036 => x"3e63417f",
  2037 => x"7f00001c",
  2038 => x"4149497f",
  2039 => x"7f000041",
  2040 => x"0109097f",
  2041 => x"3e000001",
  2042 => x"7b49417f",
  2043 => x"7f00007a",
  2044 => x"7f08087f",
  2045 => x"0000007f",
  2046 => x"417f7f41",
  2047 => x"20000000",
  2048 => x"7f404060",
  2049 => x"7f7f003f",
  2050 => x"63361c08",
  2051 => x"7f000041",
  2052 => x"4040407f",
  2053 => x"7f7f0040",
  2054 => x"7f060c06",
  2055 => x"7f7f007f",
  2056 => x"7f180c06",
  2057 => x"3e00007f",
  2058 => x"7f41417f",
  2059 => x"7f00003e",
  2060 => x"0f09097f",
  2061 => x"7f3e0006",
  2062 => x"7e7f6141",
  2063 => x"7f000040",
  2064 => x"7f19097f",
  2065 => x"26000066",
  2066 => x"7b594d6f",
  2067 => x"01000032",
  2068 => x"017f7f01",
  2069 => x"3f000001",
  2070 => x"7f40407f",
  2071 => x"0f00003f",
  2072 => x"3f70703f",
  2073 => x"7f7f000f",
  2074 => x"7f301830",
  2075 => x"6341007f",
  2076 => x"361c1c36",
  2077 => x"03014163",
  2078 => x"067c7c06",
  2079 => x"71610103",
  2080 => x"43474d59",
  2081 => x"00000041",
  2082 => x"41417f7f",
  2083 => x"03010000",
  2084 => x"30180c06",
  2085 => x"00004060",
  2086 => x"7f7f4141",
  2087 => x"0c080000",
  2088 => x"0c060306",
  2089 => x"80800008",
  2090 => x"80808080",
  2091 => x"00000080",
  2092 => x"04070300",
  2093 => x"20000000",
  2094 => x"7c545474",
  2095 => x"7f000078",
  2096 => x"7c44447f",
  2097 => x"38000038",
  2098 => x"4444447c",
  2099 => x"38000000",
  2100 => x"7f44447c",
  2101 => x"3800007f",
  2102 => x"5c54547c",
  2103 => x"04000018",
  2104 => x"05057f7e",
  2105 => x"18000000",
  2106 => x"fca4a4bc",
  2107 => x"7f00007c",
  2108 => x"7c04047f",
  2109 => x"00000078",
  2110 => x"407d3d00",
  2111 => x"80000000",
  2112 => x"7dfd8080",
  2113 => x"7f000000",
  2114 => x"6c38107f",
  2115 => x"00000044",
  2116 => x"407f3f00",
  2117 => x"7c7c0000",
  2118 => x"7c0c180c",
  2119 => x"7c000078",
  2120 => x"7c04047c",
  2121 => x"38000078",
  2122 => x"7c44447c",
  2123 => x"fc000038",
  2124 => x"3c2424fc",
  2125 => x"18000018",
  2126 => x"fc24243c",
  2127 => x"7c0000fc",
  2128 => x"0c04047c",
  2129 => x"48000008",
  2130 => x"7454545c",
  2131 => x"04000020",
  2132 => x"44447f3f",
  2133 => x"3c000000",
  2134 => x"7c40407c",
  2135 => x"1c00007c",
  2136 => x"3c60603c",
  2137 => x"7c3c001c",
  2138 => x"7c603060",
  2139 => x"6c44003c",
  2140 => x"6c381038",
  2141 => x"1c000044",
  2142 => x"3c60e0bc",
  2143 => x"4400001c",
  2144 => x"4c5c7464",
  2145 => x"08000044",
  2146 => x"41773e08",
  2147 => x"00000041",
  2148 => x"007f7f00",
  2149 => x"41000000",
  2150 => x"083e7741",
  2151 => x"01020008",
  2152 => x"02020301",
  2153 => x"7f7f0001",
  2154 => x"7f7f7f7f",
  2155 => x"0808007f",
  2156 => x"3e3e1c1c",
  2157 => x"7f7f7f7f",
  2158 => x"1c1c3e3e",
  2159 => x"10000808",
  2160 => x"187c7c18",
  2161 => x"10000010",
  2162 => x"307c7c30",
  2163 => x"30100010",
  2164 => x"1e786060",
  2165 => x"66420006",
  2166 => x"663c183c",
  2167 => x"38780042",
  2168 => x"6cc6c26a",
  2169 => x"00600038",
  2170 => x"00006000",
  2171 => x"5e0e0060",
  2172 => x"0e5d5c5b",
  2173 => x"c24c711e",
  2174 => x"4bbff6eb",
  2175 => x"48faebc2",
  2176 => x"f62778c0",
  2177 => x"bf00002a",
  2178 => x"9949bf97",
  2179 => x"87c8c102",
  2180 => x"ebc21ec0",
  2181 => x"744dbffa",
  2182 => x"87c702ad",
  2183 => x"c048a6c4",
  2184 => x"c487c578",
  2185 => x"78c148a6",
  2186 => x"751e66c4",
  2187 => x"87c4ed49",
  2188 => x"e0c086c8",
  2189 => x"87f5ee49",
  2190 => x"6a4aa3c4",
  2191 => x"87f7ef49",
  2192 => x"c287cdf0",
  2193 => x"48bffaeb",
  2194 => x"ebc280c1",
  2195 => x"83cc58fe",
  2196 => x"99496b97",
  2197 => x"87f8fe05",
  2198 => x"bffaebc2",
  2199 => x"adb7c84d",
  2200 => x"c087d903",
  2201 => x"ebc21e1e",
  2202 => x"ec49bffa",
  2203 => x"86c887c6",
  2204 => x"c187ddef",
  2205 => x"adb7c885",
  2206 => x"87e7ff04",
  2207 => x"264d2626",
  2208 => x"264b264c",
  2209 => x"4a711e4f",
  2210 => x"5afaebc2",
  2211 => x"bffeebc2",
  2212 => x"87dafd49",
  2213 => x"bffaebc2",
  2214 => x"c289c149",
  2215 => x"7159c2ec",
  2216 => x"2687cbfd",
  2217 => x"c0c11e4f",
  2218 => x"87d8ea49",
  2219 => x"48ebd6c2",
  2220 => x"4f2678c0",
  2221 => x"5c5b5e0e",
  2222 => x"86f40e5d",
  2223 => x"c048a6c8",
  2224 => x"7ebfec78",
  2225 => x"ebc280fc",
  2226 => x"c278bff6",
  2227 => x"4dbfc2ec",
  2228 => x"c74cbfe8",
  2229 => x"87f7e549",
  2230 => x"99c24970",
  2231 => x"c287cf05",
  2232 => x"49bfe3d6",
  2233 => x"996eb9ff",
  2234 => x"c00299c1",
  2235 => x"49c787ee",
  2236 => x"7087dce5",
  2237 => x"87cd0298",
  2238 => x"c787cae1",
  2239 => x"87cfe549",
  2240 => x"f3059870",
  2241 => x"ebd6c287",
  2242 => x"bac14abf",
  2243 => x"5aefd6c2",
  2244 => x"49a2c0c1",
  2245 => x"c887ede8",
  2246 => x"78c148a6",
  2247 => x"48e3d6c2",
  2248 => x"d6c2786e",
  2249 => x"c105bfeb",
  2250 => x"a6c487da",
  2251 => x"c0c0c848",
  2252 => x"efd6c278",
  2253 => x"bf976e7e",
  2254 => x"c1486e49",
  2255 => x"58a6c480",
  2256 => x"87cbe471",
  2257 => x"c3029870",
  2258 => x"b466c487",
  2259 => x"c14866c4",
  2260 => x"a6c828b7",
  2261 => x"05987058",
  2262 => x"7487daff",
  2263 => x"99ffc349",
  2264 => x"49c01e71",
  2265 => x"7487d0e6",
  2266 => x"29b7c849",
  2267 => x"49c11e71",
  2268 => x"c887c4e6",
  2269 => x"49fdc386",
  2270 => x"c387d4e3",
  2271 => x"cee349fa",
  2272 => x"87cac887",
  2273 => x"ffc34974",
  2274 => x"2cb7c899",
  2275 => x"9c74b471",
  2276 => x"ff87dd02",
  2277 => x"6e7ebfc8",
  2278 => x"e7d6c249",
  2279 => x"c0c289bf",
  2280 => x"87c403a9",
  2281 => x"87ce4cc0",
  2282 => x"48e7d6c2",
  2283 => x"87c6786e",
  2284 => x"48e7d6c2",
  2285 => x"497478c0",
  2286 => x"ce0599c8",
  2287 => x"49f5c387",
  2288 => x"7087cce2",
  2289 => x"0299c249",
  2290 => x"c287edc0",
  2291 => x"02bffeeb",
  2292 => x"c14887c9",
  2293 => x"c2ecc288",
  2294 => x"c287d858",
  2295 => x"49bffaeb",
  2296 => x"66c491cc",
  2297 => x"7ea1c881",
  2298 => x"c002bf6e",
  2299 => x"ff4b87c5",
  2300 => x"c80f7349",
  2301 => x"78c148a6",
  2302 => x"99c44974",
  2303 => x"c387ce05",
  2304 => x"cae149f2",
  2305 => x"c2497087",
  2306 => x"fdc00299",
  2307 => x"48a6c887",
  2308 => x"bffaebc2",
  2309 => x"4966c878",
  2310 => x"ebc289c1",
  2311 => x"6e7ebffe",
  2312 => x"c006a9b7",
  2313 => x"c14887c9",
  2314 => x"c2ecc280",
  2315 => x"c887d658",
  2316 => x"91cc4966",
  2317 => x"c88166c4",
  2318 => x"bf6e7ea1",
  2319 => x"87c5c002",
  2320 => x"7349fe4b",
  2321 => x"48a6c80f",
  2322 => x"fdc378c1",
  2323 => x"fedfff49",
  2324 => x"c2497087",
  2325 => x"eec00299",
  2326 => x"feebc287",
  2327 => x"c9c002bf",
  2328 => x"feebc287",
  2329 => x"c078c048",
  2330 => x"ebc287d8",
  2331 => x"cc49bffa",
  2332 => x"8166c491",
  2333 => x"6e7ea1c8",
  2334 => x"c5c002bf",
  2335 => x"49fd4b87",
  2336 => x"a6c80f73",
  2337 => x"c378c148",
  2338 => x"dfff49fa",
  2339 => x"497087c1",
  2340 => x"c10299c2",
  2341 => x"a6c887c0",
  2342 => x"faebc248",
  2343 => x"66c878bf",
  2344 => x"c488c148",
  2345 => x"ebc258a6",
  2346 => x"6e48bffe",
  2347 => x"c003a8b7",
  2348 => x"ebc287c9",
  2349 => x"786e48fe",
  2350 => x"c887d6c0",
  2351 => x"91cc4966",
  2352 => x"c88166c4",
  2353 => x"bf6e7ea1",
  2354 => x"87c5c002",
  2355 => x"7349fc4b",
  2356 => x"48a6c80f",
  2357 => x"ebc278c1",
  2358 => x"c04abffe",
  2359 => x"c006aab7",
  2360 => x"8ac187c9",
  2361 => x"01aab7c0",
  2362 => x"7487f7ff",
  2363 => x"99f0c349",
  2364 => x"87cfc005",
  2365 => x"ff49dac1",
  2366 => x"7087d4dd",
  2367 => x"0299c249",
  2368 => x"c287cec1",
  2369 => x"7ebff6eb",
  2370 => x"c248a6c4",
  2371 => x"78bffeeb",
  2372 => x"484a66c4",
  2373 => x"06a8b7c0",
  2374 => x"6e87d0c0",
  2375 => x"c480cc48",
  2376 => x"8ac158a6",
  2377 => x"01aab7c0",
  2378 => x"6e87f0ff",
  2379 => x"c24bbf97",
  2380 => x"d1c0028b",
  2381 => x"c0058b87",
  2382 => x"4a6e87d7",
  2383 => x"496a82c8",
  2384 => x"c087c2f5",
  2385 => x"4b6e87cb",
  2386 => x"4b6b83c8",
  2387 => x"734966c4",
  2388 => x"029d750f",
  2389 => x"6d87e9c0",
  2390 => x"87e4c002",
  2391 => x"dbff496d",
  2392 => x"497087ed",
  2393 => x"c00299c1",
  2394 => x"a5c487cb",
  2395 => x"feebc24b",
  2396 => x"4b6b49bf",
  2397 => x"0285c80f",
  2398 => x"6d87c5c0",
  2399 => x"87dcff05",
  2400 => x"c00266c8",
  2401 => x"ebc287c8",
  2402 => x"f149bffe",
  2403 => x"8ef487e0",
  2404 => x"5887eaf3",
  2405 => x"1d141112",
  2406 => x"5a231c1b",
  2407 => x"f5949159",
  2408 => x"00f4ebf2",
  2409 => x"00000000",
  2410 => x"00000000",
  2411 => x"58000000",
  2412 => x"1d111412",
  2413 => x"5a231c1b",
  2414 => x"f5919459",
  2415 => x"00f4ebf2",
  2416 => x"000025c4",
  2417 => x"4f545541",
  2418 => x"544f4f42",
  2419 => x"0053454e",
  2420 => x"000019c4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
