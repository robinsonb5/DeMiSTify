
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c8",x"ec",x"c2",x"87"),
    12 => (x"86",x"c0",x"c4",x"4e"),
    13 => (x"49",x"c8",x"ec",x"c2"),
    14 => (x"48",x"d4",x"d7",x"c2"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"d4",x"d7",x"c2",x"87"),
    21 => (x"d0",x"d7",x"c2",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"e1",x"c1",x"87",x"f7"),
    25 => (x"d7",x"c2",x"87",x"c1"),
    26 => (x"d7",x"c2",x"4d",x"d4"),
    27 => (x"ad",x"74",x"4c",x"d4"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"5c",x"5b",x"5e",x"0e"),
    32 => (x"c0",x"4b",x"71",x"0e"),
    33 => (x"9a",x"4a",x"13",x"4c"),
    34 => (x"72",x"87",x"cd",x"02"),
    35 => (x"87",x"e0",x"c0",x"49"),
    36 => (x"4a",x"13",x"84",x"c1"),
    37 => (x"87",x"f3",x"05",x"9a"),
    38 => (x"4c",x"26",x"48",x"74"),
    39 => (x"4f",x"26",x"4b",x"26"),
    40 => (x"81",x"48",x"73",x"1e"),
    41 => (x"c5",x"02",x"a9",x"73"),
    42 => (x"05",x"53",x"12",x"87"),
    43 => (x"4f",x"26",x"87",x"f6"),
    44 => (x"c0",x"ff",x"1e",x"1e"),
    45 => (x"c4",x"48",x"6a",x"4a"),
    46 => (x"a6",x"c4",x"98",x"c0"),
    47 => (x"02",x"98",x"70",x"58"),
    48 => (x"7a",x"71",x"87",x"f3"),
    49 => (x"4f",x"26",x"26",x"48"),
    50 => (x"ff",x"1e",x"73",x"1e"),
    51 => (x"ff",x"c3",x"4b",x"d4"),
    52 => (x"c3",x"4a",x"6b",x"7b"),
    53 => (x"49",x"6b",x"7b",x"ff"),
    54 => (x"b1",x"72",x"32",x"c8"),
    55 => (x"6b",x"7b",x"ff",x"c3"),
    56 => (x"71",x"31",x"c8",x"4a"),
    57 => (x"7b",x"ff",x"c3",x"b2"),
    58 => (x"32",x"c8",x"49",x"6b"),
    59 => (x"48",x"71",x"b1",x"72"),
    60 => (x"4d",x"26",x"87",x"c4"),
    61 => (x"4b",x"26",x"4c",x"26"),
    62 => (x"5e",x"0e",x"4f",x"26"),
    63 => (x"0e",x"5d",x"5c",x"5b"),
    64 => (x"d4",x"ff",x"4a",x"71"),
    65 => (x"c3",x"48",x"72",x"4c"),
    66 => (x"7c",x"70",x"98",x"ff"),
    67 => (x"bf",x"d4",x"d7",x"c2"),
    68 => (x"d0",x"87",x"c8",x"05"),
    69 => (x"30",x"c9",x"48",x"66"),
    70 => (x"d0",x"58",x"a6",x"d4"),
    71 => (x"29",x"d8",x"49",x"66"),
    72 => (x"ff",x"c3",x"48",x"71"),
    73 => (x"d0",x"7c",x"70",x"98"),
    74 => (x"29",x"d0",x"49",x"66"),
    75 => (x"ff",x"c3",x"48",x"71"),
    76 => (x"d0",x"7c",x"70",x"98"),
    77 => (x"29",x"c8",x"49",x"66"),
    78 => (x"ff",x"c3",x"48",x"71"),
    79 => (x"d0",x"7c",x"70",x"98"),
    80 => (x"ff",x"c3",x"48",x"66"),
    81 => (x"72",x"7c",x"70",x"98"),
    82 => (x"71",x"29",x"d0",x"49"),
    83 => (x"98",x"ff",x"c3",x"48"),
    84 => (x"4b",x"6c",x"7c",x"70"),
    85 => (x"4d",x"ff",x"f0",x"c9"),
    86 => (x"05",x"ab",x"ff",x"c3"),
    87 => (x"ff",x"c3",x"87",x"d0"),
    88 => (x"c1",x"4b",x"6c",x"7c"),
    89 => (x"87",x"c6",x"02",x"8d"),
    90 => (x"02",x"ab",x"ff",x"c3"),
    91 => (x"48",x"73",x"87",x"f0"),
    92 => (x"1e",x"87",x"ff",x"fd"),
    93 => (x"d4",x"ff",x"49",x"c0"),
    94 => (x"78",x"ff",x"c3",x"48"),
    95 => (x"c8",x"c3",x"81",x"c1"),
    96 => (x"f1",x"04",x"a9",x"b7"),
    97 => (x"1e",x"4f",x"26",x"87"),
    98 => (x"87",x"e7",x"1e",x"73"),
    99 => (x"4b",x"df",x"f8",x"c4"),
   100 => (x"ff",x"c0",x"1e",x"c0"),
   101 => (x"49",x"f7",x"c1",x"f0"),
   102 => (x"c4",x"87",x"df",x"fd"),
   103 => (x"05",x"a8",x"c1",x"86"),
   104 => (x"ff",x"87",x"ea",x"c0"),
   105 => (x"ff",x"c3",x"48",x"d4"),
   106 => (x"c0",x"c0",x"c1",x"78"),
   107 => (x"1e",x"c0",x"c0",x"c0"),
   108 => (x"c1",x"f0",x"e1",x"c0"),
   109 => (x"c1",x"fd",x"49",x"e9"),
   110 => (x"70",x"86",x"c4",x"87"),
   111 => (x"87",x"ca",x"05",x"98"),
   112 => (x"c3",x"48",x"d4",x"ff"),
   113 => (x"48",x"c1",x"78",x"ff"),
   114 => (x"e6",x"fe",x"87",x"cb"),
   115 => (x"05",x"8b",x"c1",x"87"),
   116 => (x"c0",x"87",x"fd",x"fe"),
   117 => (x"87",x"de",x"fc",x"48"),
   118 => (x"ff",x"1e",x"73",x"1e"),
   119 => (x"ff",x"c3",x"48",x"d4"),
   120 => (x"49",x"d3",x"c8",x"78"),
   121 => (x"d3",x"87",x"d5",x"fa"),
   122 => (x"c0",x"1e",x"c0",x"4b"),
   123 => (x"c1",x"c1",x"f0",x"ff"),
   124 => (x"87",x"c6",x"fc",x"49"),
   125 => (x"98",x"70",x"86",x"c4"),
   126 => (x"ff",x"87",x"ca",x"05"),
   127 => (x"ff",x"c3",x"48",x"d4"),
   128 => (x"cb",x"48",x"c1",x"78"),
   129 => (x"87",x"eb",x"fd",x"87"),
   130 => (x"ff",x"05",x"8b",x"c1"),
   131 => (x"48",x"c0",x"87",x"db"),
   132 => (x"43",x"87",x"e3",x"fb"),
   133 => (x"53",x"00",x"44",x"4d"),
   134 => (x"20",x"43",x"48",x"44"),
   135 => (x"6c",x"69",x"61",x"66"),
   136 => (x"49",x"00",x"0a",x"21"),
   137 => (x"00",x"52",x"52",x"45"),
   138 => (x"00",x"49",x"50",x"53"),
   139 => (x"74",x"69",x"72",x"57"),
   140 => (x"61",x"66",x"20",x"65"),
   141 => (x"64",x"65",x"6c",x"69"),
   142 => (x"5e",x"0e",x"00",x"0a"),
   143 => (x"ff",x"0e",x"5c",x"5b"),
   144 => (x"ee",x"fc",x"4c",x"d4"),
   145 => (x"1e",x"ea",x"c6",x"87"),
   146 => (x"c1",x"f0",x"e1",x"c0"),
   147 => (x"e9",x"fa",x"49",x"c8"),
   148 => (x"c1",x"86",x"c4",x"87"),
   149 => (x"87",x"c8",x"02",x"a8"),
   150 => (x"c0",x"87",x"fd",x"fd"),
   151 => (x"87",x"e8",x"c1",x"48"),
   152 => (x"70",x"87",x"e5",x"f9"),
   153 => (x"ff",x"ff",x"cf",x"49"),
   154 => (x"a9",x"ea",x"c6",x"99"),
   155 => (x"fd",x"87",x"c8",x"02"),
   156 => (x"48",x"c0",x"87",x"e6"),
   157 => (x"c3",x"87",x"d1",x"c1"),
   158 => (x"f1",x"c0",x"7c",x"ff"),
   159 => (x"87",x"c7",x"fc",x"4b"),
   160 => (x"c0",x"02",x"98",x"70"),
   161 => (x"1e",x"c0",x"87",x"eb"),
   162 => (x"c1",x"f0",x"ff",x"c0"),
   163 => (x"e9",x"f9",x"49",x"fa"),
   164 => (x"70",x"86",x"c4",x"87"),
   165 => (x"87",x"d9",x"05",x"98"),
   166 => (x"6c",x"7c",x"ff",x"c3"),
   167 => (x"7c",x"ff",x"c3",x"49"),
   168 => (x"c1",x"7c",x"7c",x"7c"),
   169 => (x"c4",x"02",x"99",x"c0"),
   170 => (x"db",x"48",x"c1",x"87"),
   171 => (x"d7",x"48",x"c0",x"87"),
   172 => (x"05",x"ab",x"c2",x"87"),
   173 => (x"d7",x"c8",x"87",x"ca"),
   174 => (x"87",x"c0",x"f7",x"49"),
   175 => (x"87",x"c8",x"48",x"c0"),
   176 => (x"fe",x"05",x"8b",x"c1"),
   177 => (x"48",x"c0",x"87",x"f7"),
   178 => (x"0e",x"87",x"e9",x"f8"),
   179 => (x"5d",x"5c",x"5b",x"5e"),
   180 => (x"d0",x"ff",x"1e",x"0e"),
   181 => (x"c0",x"c0",x"c8",x"4d"),
   182 => (x"d4",x"d7",x"c2",x"4b"),
   183 => (x"c8",x"78",x"c1",x"48"),
   184 => (x"d7",x"f6",x"49",x"e8"),
   185 => (x"6d",x"4c",x"c7",x"87"),
   186 => (x"c4",x"98",x"73",x"48"),
   187 => (x"98",x"70",x"58",x"a6"),
   188 => (x"6d",x"87",x"cc",x"02"),
   189 => (x"c4",x"98",x"73",x"48"),
   190 => (x"98",x"70",x"58",x"a6"),
   191 => (x"c2",x"87",x"f4",x"05"),
   192 => (x"87",x"ef",x"f9",x"7d"),
   193 => (x"98",x"73",x"48",x"6d"),
   194 => (x"70",x"58",x"a6",x"c4"),
   195 => (x"87",x"cc",x"02",x"98"),
   196 => (x"98",x"73",x"48",x"6d"),
   197 => (x"70",x"58",x"a6",x"c4"),
   198 => (x"87",x"f4",x"05",x"98"),
   199 => (x"1e",x"c0",x"7d",x"c3"),
   200 => (x"c1",x"d0",x"e5",x"c0"),
   201 => (x"d1",x"f7",x"49",x"c0"),
   202 => (x"c1",x"86",x"c4",x"87"),
   203 => (x"87",x"c1",x"05",x"a8"),
   204 => (x"05",x"ac",x"c2",x"4c"),
   205 => (x"e3",x"c8",x"87",x"cb"),
   206 => (x"87",x"c0",x"f5",x"49"),
   207 => (x"ce",x"c1",x"48",x"c0"),
   208 => (x"05",x"8c",x"c1",x"87"),
   209 => (x"fb",x"87",x"e0",x"fe"),
   210 => (x"d7",x"c2",x"87",x"f0"),
   211 => (x"98",x"70",x"58",x"d8"),
   212 => (x"c1",x"87",x"cd",x"05"),
   213 => (x"f0",x"ff",x"c0",x"1e"),
   214 => (x"f6",x"49",x"d0",x"c1"),
   215 => (x"86",x"c4",x"87",x"dc"),
   216 => (x"c3",x"48",x"d4",x"ff"),
   217 => (x"dd",x"c5",x"78",x"ff"),
   218 => (x"dc",x"d7",x"c2",x"87"),
   219 => (x"73",x"48",x"6d",x"58"),
   220 => (x"58",x"a6",x"c4",x"98"),
   221 => (x"cc",x"02",x"98",x"70"),
   222 => (x"73",x"48",x"6d",x"87"),
   223 => (x"58",x"a6",x"c4",x"98"),
   224 => (x"f4",x"05",x"98",x"70"),
   225 => (x"ff",x"7d",x"c2",x"87"),
   226 => (x"ff",x"c3",x"48",x"d4"),
   227 => (x"26",x"48",x"c1",x"78"),
   228 => (x"0e",x"87",x"df",x"f5"),
   229 => (x"5d",x"5c",x"5b",x"5e"),
   230 => (x"c0",x"c8",x"1e",x"0e"),
   231 => (x"4c",x"c0",x"4b",x"c0"),
   232 => (x"df",x"cd",x"ee",x"c5"),
   233 => (x"5c",x"a6",x"c4",x"4a"),
   234 => (x"c3",x"4c",x"d4",x"ff"),
   235 => (x"48",x"6c",x"7c",x"ff"),
   236 => (x"05",x"a8",x"fe",x"c3"),
   237 => (x"71",x"87",x"c0",x"c2"),
   238 => (x"e2",x"c0",x"05",x"99"),
   239 => (x"bf",x"d0",x"ff",x"87"),
   240 => (x"c4",x"98",x"73",x"48"),
   241 => (x"98",x"70",x"58",x"a6"),
   242 => (x"ff",x"87",x"ce",x"02"),
   243 => (x"73",x"48",x"bf",x"d0"),
   244 => (x"58",x"a6",x"c4",x"98"),
   245 => (x"f2",x"05",x"98",x"70"),
   246 => (x"48",x"d0",x"ff",x"87"),
   247 => (x"d4",x"78",x"d1",x"c4"),
   248 => (x"b7",x"c0",x"48",x"66"),
   249 => (x"e0",x"c0",x"06",x"a8"),
   250 => (x"7c",x"ff",x"c3",x"87"),
   251 => (x"99",x"71",x"4a",x"6c"),
   252 => (x"71",x"87",x"c7",x"02"),
   253 => (x"0a",x"7a",x"97",x"0a"),
   254 => (x"66",x"d4",x"81",x"c1"),
   255 => (x"d8",x"88",x"c1",x"48"),
   256 => (x"b7",x"c0",x"58",x"a6"),
   257 => (x"e0",x"ff",x"01",x"a8"),
   258 => (x"7c",x"ff",x"c3",x"87"),
   259 => (x"05",x"99",x"71",x"7c"),
   260 => (x"ff",x"87",x"e1",x"c0"),
   261 => (x"73",x"48",x"bf",x"d0"),
   262 => (x"58",x"a6",x"c4",x"98"),
   263 => (x"ce",x"02",x"98",x"70"),
   264 => (x"bf",x"d0",x"ff",x"87"),
   265 => (x"c4",x"98",x"73",x"48"),
   266 => (x"98",x"70",x"58",x"a6"),
   267 => (x"ff",x"87",x"f2",x"05"),
   268 => (x"78",x"d0",x"48",x"d0"),
   269 => (x"c1",x"7e",x"4a",x"c1"),
   270 => (x"ee",x"fd",x"05",x"8a"),
   271 => (x"26",x"48",x"6e",x"87"),
   272 => (x"0e",x"87",x"ef",x"f2"),
   273 => (x"0e",x"5c",x"5b",x"5e"),
   274 => (x"c8",x"4a",x"71",x"1e"),
   275 => (x"c0",x"4b",x"c0",x"c0"),
   276 => (x"48",x"d4",x"ff",x"4c"),
   277 => (x"ff",x"78",x"ff",x"c3"),
   278 => (x"73",x"48",x"bf",x"d0"),
   279 => (x"58",x"a6",x"c4",x"98"),
   280 => (x"ce",x"02",x"98",x"70"),
   281 => (x"bf",x"d0",x"ff",x"87"),
   282 => (x"c4",x"98",x"73",x"48"),
   283 => (x"98",x"70",x"58",x"a6"),
   284 => (x"ff",x"87",x"f2",x"05"),
   285 => (x"c3",x"c4",x"48",x"d0"),
   286 => (x"48",x"d4",x"ff",x"78"),
   287 => (x"72",x"78",x"ff",x"c3"),
   288 => (x"f0",x"ff",x"c0",x"1e"),
   289 => (x"f1",x"49",x"d1",x"c1"),
   290 => (x"86",x"c4",x"87",x"f0"),
   291 => (x"c0",x"05",x"98",x"70"),
   292 => (x"c0",x"c8",x"87",x"ee"),
   293 => (x"49",x"66",x"d4",x"1e"),
   294 => (x"c4",x"87",x"f8",x"fb"),
   295 => (x"ff",x"4c",x"70",x"86"),
   296 => (x"73",x"48",x"bf",x"d0"),
   297 => (x"58",x"a6",x"c4",x"98"),
   298 => (x"ce",x"02",x"98",x"70"),
   299 => (x"bf",x"d0",x"ff",x"87"),
   300 => (x"c4",x"98",x"73",x"48"),
   301 => (x"98",x"70",x"58",x"a6"),
   302 => (x"ff",x"87",x"f2",x"05"),
   303 => (x"78",x"c2",x"48",x"d0"),
   304 => (x"f0",x"26",x"48",x"74"),
   305 => (x"5e",x"0e",x"87",x"ee"),
   306 => (x"0e",x"5d",x"5c",x"5b"),
   307 => (x"ff",x"c0",x"1e",x"c0"),
   308 => (x"49",x"c9",x"c1",x"f0"),
   309 => (x"d2",x"87",x"e3",x"f0"),
   310 => (x"e2",x"d7",x"c2",x"1e"),
   311 => (x"87",x"f3",x"fa",x"49"),
   312 => (x"4c",x"c0",x"86",x"c8"),
   313 => (x"b7",x"d2",x"84",x"c1"),
   314 => (x"87",x"f8",x"04",x"ac"),
   315 => (x"97",x"e2",x"d7",x"c2"),
   316 => (x"c0",x"c3",x"49",x"bf"),
   317 => (x"a9",x"c0",x"c1",x"99"),
   318 => (x"87",x"e7",x"c0",x"05"),
   319 => (x"97",x"e9",x"d7",x"c2"),
   320 => (x"31",x"d0",x"49",x"bf"),
   321 => (x"97",x"ea",x"d7",x"c2"),
   322 => (x"32",x"c8",x"4a",x"bf"),
   323 => (x"d7",x"c2",x"b1",x"72"),
   324 => (x"4a",x"bf",x"97",x"eb"),
   325 => (x"cf",x"4c",x"71",x"b1"),
   326 => (x"9c",x"ff",x"ff",x"ff"),
   327 => (x"34",x"ca",x"84",x"c1"),
   328 => (x"c2",x"87",x"e7",x"c1"),
   329 => (x"bf",x"97",x"eb",x"d7"),
   330 => (x"c6",x"31",x"c1",x"49"),
   331 => (x"ec",x"d7",x"c2",x"99"),
   332 => (x"c7",x"4a",x"bf",x"97"),
   333 => (x"b1",x"72",x"2a",x"b7"),
   334 => (x"97",x"e7",x"d7",x"c2"),
   335 => (x"cf",x"4d",x"4a",x"bf"),
   336 => (x"e8",x"d7",x"c2",x"9d"),
   337 => (x"c3",x"4a",x"bf",x"97"),
   338 => (x"c2",x"32",x"ca",x"9a"),
   339 => (x"bf",x"97",x"e9",x"d7"),
   340 => (x"73",x"33",x"c2",x"4b"),
   341 => (x"ea",x"d7",x"c2",x"b2"),
   342 => (x"c3",x"4b",x"bf",x"97"),
   343 => (x"b7",x"c6",x"9b",x"c0"),
   344 => (x"c2",x"b2",x"73",x"2b"),
   345 => (x"71",x"48",x"c1",x"81"),
   346 => (x"c1",x"49",x"70",x"30"),
   347 => (x"70",x"30",x"75",x"48"),
   348 => (x"c1",x"4c",x"72",x"4d"),
   349 => (x"c8",x"94",x"71",x"84"),
   350 => (x"06",x"ad",x"b7",x"c0"),
   351 => (x"34",x"c1",x"87",x"cc"),
   352 => (x"c0",x"c8",x"2d",x"b7"),
   353 => (x"ff",x"01",x"ad",x"b7"),
   354 => (x"48",x"74",x"87",x"f4"),
   355 => (x"0e",x"87",x"e3",x"ed"),
   356 => (x"0e",x"5c",x"5b",x"5e"),
   357 => (x"4c",x"c0",x"4b",x"71"),
   358 => (x"c0",x"48",x"66",x"d0"),
   359 => (x"c0",x"06",x"a8",x"b7"),
   360 => (x"4a",x"13",x"87",x"e3"),
   361 => (x"bf",x"97",x"66",x"cc"),
   362 => (x"48",x"66",x"cc",x"49"),
   363 => (x"a6",x"d0",x"80",x"c1"),
   364 => (x"aa",x"b7",x"71",x"58"),
   365 => (x"c1",x"87",x"c4",x"02"),
   366 => (x"c1",x"87",x"cc",x"48"),
   367 => (x"b7",x"66",x"d0",x"84"),
   368 => (x"dd",x"ff",x"04",x"ac"),
   369 => (x"c2",x"48",x"c0",x"87"),
   370 => (x"26",x"4d",x"26",x"87"),
   371 => (x"26",x"4b",x"26",x"4c"),
   372 => (x"5b",x"5e",x"0e",x"4f"),
   373 => (x"c2",x"0e",x"5d",x"5c"),
   374 => (x"c0",x"48",x"c8",x"e0"),
   375 => (x"c0",x"d8",x"c2",x"78"),
   376 => (x"f9",x"49",x"c0",x"1e"),
   377 => (x"86",x"c4",x"87",x"dd"),
   378 => (x"c5",x"05",x"98",x"70"),
   379 => (x"c8",x"48",x"c0",x"87"),
   380 => (x"4b",x"c0",x"87",x"ef"),
   381 => (x"48",x"c0",x"e5",x"c2"),
   382 => (x"1e",x"c8",x"78",x"c1"),
   383 => (x"1e",x"ed",x"e0",x"c0"),
   384 => (x"49",x"f6",x"d8",x"c2"),
   385 => (x"c8",x"87",x"c8",x"fe"),
   386 => (x"05",x"98",x"70",x"86"),
   387 => (x"e5",x"c2",x"87",x"c6"),
   388 => (x"78",x"c0",x"48",x"c0"),
   389 => (x"e0",x"c0",x"1e",x"c8"),
   390 => (x"d9",x"c2",x"1e",x"f6"),
   391 => (x"ee",x"fd",x"49",x"d2"),
   392 => (x"70",x"86",x"c8",x"87"),
   393 => (x"87",x"c6",x"05",x"98"),
   394 => (x"48",x"c0",x"e5",x"c2"),
   395 => (x"e5",x"c2",x"78",x"c0"),
   396 => (x"c0",x"02",x"bf",x"c0"),
   397 => (x"df",x"c2",x"87",x"fa"),
   398 => (x"c2",x"4b",x"bf",x"c6"),
   399 => (x"bf",x"9f",x"fe",x"df"),
   400 => (x"ea",x"d6",x"c5",x"4a"),
   401 => (x"87",x"c7",x"05",x"aa"),
   402 => (x"bf",x"c6",x"df",x"c2"),
   403 => (x"ca",x"87",x"cc",x"4b"),
   404 => (x"02",x"aa",x"d5",x"e9"),
   405 => (x"48",x"c0",x"87",x"c5"),
   406 => (x"c2",x"87",x"c6",x"c7"),
   407 => (x"73",x"1e",x"c0",x"d8"),
   408 => (x"87",x"df",x"f7",x"49"),
   409 => (x"98",x"70",x"86",x"c4"),
   410 => (x"c0",x"87",x"c5",x"05"),
   411 => (x"87",x"f1",x"c6",x"48"),
   412 => (x"e0",x"c0",x"1e",x"c8"),
   413 => (x"d9",x"c2",x"1e",x"ff"),
   414 => (x"d2",x"fc",x"49",x"d2"),
   415 => (x"70",x"86",x"c8",x"87"),
   416 => (x"87",x"c8",x"05",x"98"),
   417 => (x"48",x"c8",x"e0",x"c2"),
   418 => (x"87",x"da",x"78",x"c1"),
   419 => (x"e1",x"c0",x"1e",x"c8"),
   420 => (x"d8",x"c2",x"1e",x"c8"),
   421 => (x"f6",x"fb",x"49",x"f6"),
   422 => (x"70",x"86",x"c8",x"87"),
   423 => (x"c5",x"c0",x"02",x"98"),
   424 => (x"c5",x"48",x"c0",x"87"),
   425 => (x"df",x"c2",x"87",x"fb"),
   426 => (x"49",x"bf",x"97",x"fe"),
   427 => (x"05",x"a9",x"d5",x"c1"),
   428 => (x"c2",x"87",x"cd",x"c0"),
   429 => (x"bf",x"97",x"ff",x"df"),
   430 => (x"a9",x"ea",x"c2",x"49"),
   431 => (x"87",x"c5",x"c0",x"02"),
   432 => (x"dc",x"c5",x"48",x"c0"),
   433 => (x"c0",x"d8",x"c2",x"87"),
   434 => (x"c3",x"4c",x"bf",x"97"),
   435 => (x"c0",x"02",x"ac",x"e9"),
   436 => (x"eb",x"c3",x"87",x"cc"),
   437 => (x"c5",x"c0",x"02",x"ac"),
   438 => (x"c5",x"48",x"c0",x"87"),
   439 => (x"d8",x"c2",x"87",x"c3"),
   440 => (x"49",x"bf",x"97",x"cb"),
   441 => (x"cc",x"c0",x"05",x"99"),
   442 => (x"cc",x"d8",x"c2",x"87"),
   443 => (x"c2",x"49",x"bf",x"97"),
   444 => (x"c5",x"c0",x"02",x"a9"),
   445 => (x"c4",x"48",x"c0",x"87"),
   446 => (x"d8",x"c2",x"87",x"e7"),
   447 => (x"48",x"bf",x"97",x"cd"),
   448 => (x"58",x"c4",x"e0",x"c2"),
   449 => (x"e0",x"c2",x"88",x"c1"),
   450 => (x"d8",x"c2",x"58",x"c8"),
   451 => (x"49",x"bf",x"97",x"ce"),
   452 => (x"d8",x"c2",x"81",x"73"),
   453 => (x"4a",x"bf",x"97",x"cf"),
   454 => (x"71",x"35",x"c8",x"4d"),
   455 => (x"e0",x"e4",x"c2",x"85"),
   456 => (x"d0",x"d8",x"c2",x"5d"),
   457 => (x"c2",x"48",x"bf",x"97"),
   458 => (x"c2",x"58",x"f4",x"e4"),
   459 => (x"02",x"bf",x"c8",x"e0"),
   460 => (x"c8",x"87",x"dc",x"c2"),
   461 => (x"e4",x"e0",x"c0",x"1e"),
   462 => (x"d2",x"d9",x"c2",x"1e"),
   463 => (x"87",x"cf",x"f9",x"49"),
   464 => (x"98",x"70",x"86",x"c8"),
   465 => (x"87",x"c5",x"c0",x"02"),
   466 => (x"d4",x"c3",x"48",x"c0"),
   467 => (x"c0",x"e0",x"c2",x"87"),
   468 => (x"c4",x"48",x"4a",x"bf"),
   469 => (x"d0",x"e0",x"c2",x"30"),
   470 => (x"f0",x"e4",x"c2",x"58"),
   471 => (x"e5",x"d8",x"c2",x"5a"),
   472 => (x"c8",x"49",x"bf",x"97"),
   473 => (x"e4",x"d8",x"c2",x"31"),
   474 => (x"a1",x"4b",x"bf",x"97"),
   475 => (x"e6",x"d8",x"c2",x"49"),
   476 => (x"d0",x"4b",x"bf",x"97"),
   477 => (x"49",x"a1",x"73",x"33"),
   478 => (x"97",x"e7",x"d8",x"c2"),
   479 => (x"33",x"d8",x"4b",x"bf"),
   480 => (x"c2",x"49",x"a1",x"73"),
   481 => (x"c2",x"59",x"f8",x"e4"),
   482 => (x"91",x"bf",x"f0",x"e4"),
   483 => (x"bf",x"dc",x"e4",x"c2"),
   484 => (x"e4",x"e4",x"c2",x"81"),
   485 => (x"ed",x"d8",x"c2",x"59"),
   486 => (x"c8",x"4b",x"bf",x"97"),
   487 => (x"ec",x"d8",x"c2",x"33"),
   488 => (x"a3",x"4c",x"bf",x"97"),
   489 => (x"ee",x"d8",x"c2",x"4b"),
   490 => (x"d0",x"4c",x"bf",x"97"),
   491 => (x"4b",x"a3",x"74",x"34"),
   492 => (x"97",x"ef",x"d8",x"c2"),
   493 => (x"9c",x"cf",x"4c",x"bf"),
   494 => (x"a3",x"74",x"34",x"d8"),
   495 => (x"e8",x"e4",x"c2",x"4b"),
   496 => (x"73",x"8b",x"c2",x"5b"),
   497 => (x"e8",x"e4",x"c2",x"92"),
   498 => (x"78",x"a1",x"72",x"48"),
   499 => (x"c2",x"87",x"cb",x"c1"),
   500 => (x"bf",x"97",x"d2",x"d8"),
   501 => (x"c2",x"31",x"c8",x"49"),
   502 => (x"bf",x"97",x"d1",x"d8"),
   503 => (x"c2",x"49",x"a1",x"4a"),
   504 => (x"c5",x"59",x"d0",x"e0"),
   505 => (x"81",x"ff",x"c7",x"31"),
   506 => (x"e4",x"c2",x"29",x"c9"),
   507 => (x"d8",x"c2",x"59",x"f0"),
   508 => (x"4a",x"bf",x"97",x"d7"),
   509 => (x"d8",x"c2",x"32",x"c8"),
   510 => (x"4b",x"bf",x"97",x"d6"),
   511 => (x"e4",x"c2",x"4a",x"a2"),
   512 => (x"e4",x"c2",x"5a",x"f8"),
   513 => (x"75",x"92",x"bf",x"f0"),
   514 => (x"ec",x"e4",x"c2",x"82"),
   515 => (x"e4",x"e4",x"c2",x"5a"),
   516 => (x"c2",x"78",x"c0",x"48"),
   517 => (x"72",x"48",x"e0",x"e4"),
   518 => (x"49",x"c0",x"78",x"a1"),
   519 => (x"c1",x"87",x"f7",x"c7"),
   520 => (x"87",x"e5",x"f6",x"48"),
   521 => (x"33",x"54",x"41",x"46"),
   522 => (x"20",x"20",x"20",x"32"),
   523 => (x"54",x"41",x"46",x"00"),
   524 => (x"20",x"20",x"36",x"31"),
   525 => (x"41",x"46",x"00",x"20"),
   526 => (x"20",x"32",x"33",x"54"),
   527 => (x"46",x"00",x"20",x"20"),
   528 => (x"32",x"33",x"54",x"41"),
   529 => (x"00",x"20",x"20",x"20"),
   530 => (x"31",x"54",x"41",x"46"),
   531 => (x"20",x"20",x"20",x"36"),
   532 => (x"5b",x"5e",x"0e",x"00"),
   533 => (x"71",x"0e",x"5d",x"5c"),
   534 => (x"c8",x"e0",x"c2",x"4a"),
   535 => (x"87",x"cc",x"02",x"bf"),
   536 => (x"b7",x"c7",x"4b",x"72"),
   537 => (x"c1",x"4d",x"72",x"2b"),
   538 => (x"87",x"ca",x"9d",x"ff"),
   539 => (x"b7",x"c8",x"4b",x"72"),
   540 => (x"c3",x"4d",x"72",x"2b"),
   541 => (x"d8",x"c2",x"9d",x"ff"),
   542 => (x"e4",x"c2",x"1e",x"c0"),
   543 => (x"73",x"49",x"bf",x"dc"),
   544 => (x"fe",x"ee",x"71",x"81"),
   545 => (x"70",x"86",x"c4",x"87"),
   546 => (x"87",x"c5",x"05",x"98"),
   547 => (x"e6",x"c0",x"48",x"c0"),
   548 => (x"c8",x"e0",x"c2",x"87"),
   549 => (x"87",x"d2",x"02",x"bf"),
   550 => (x"91",x"c4",x"49",x"75"),
   551 => (x"81",x"c0",x"d8",x"c2"),
   552 => (x"ff",x"cf",x"4c",x"69"),
   553 => (x"9c",x"ff",x"ff",x"ff"),
   554 => (x"49",x"75",x"87",x"cb"),
   555 => (x"d8",x"c2",x"91",x"c2"),
   556 => (x"69",x"9f",x"81",x"c0"),
   557 => (x"f4",x"48",x"74",x"4c"),
   558 => (x"5e",x"0e",x"87",x"cf"),
   559 => (x"0e",x"5d",x"5c",x"5b"),
   560 => (x"4c",x"71",x"86",x"f4"),
   561 => (x"e4",x"c2",x"4b",x"c0"),
   562 => (x"c4",x"7e",x"bf",x"f8"),
   563 => (x"e4",x"c2",x"48",x"a6"),
   564 => (x"c8",x"78",x"bf",x"fc"),
   565 => (x"78",x"c0",x"48",x"a6"),
   566 => (x"bf",x"cc",x"e0",x"c2"),
   567 => (x"06",x"a8",x"c0",x"48"),
   568 => (x"c8",x"87",x"dd",x"c2"),
   569 => (x"99",x"cf",x"49",x"66"),
   570 => (x"c2",x"87",x"d8",x"05"),
   571 => (x"c8",x"1e",x"c0",x"d8"),
   572 => (x"c1",x"48",x"49",x"66"),
   573 => (x"58",x"a6",x"cc",x"80"),
   574 => (x"c4",x"87",x"c8",x"ed"),
   575 => (x"c0",x"d8",x"c2",x"86"),
   576 => (x"c0",x"87",x"c3",x"4b"),
   577 => (x"6b",x"97",x"83",x"e0"),
   578 => (x"c1",x"02",x"9a",x"4a"),
   579 => (x"e5",x"c3",x"87",x"e1"),
   580 => (x"da",x"c1",x"02",x"aa"),
   581 => (x"49",x"a3",x"cb",x"87"),
   582 => (x"d8",x"49",x"69",x"97"),
   583 => (x"ce",x"c1",x"05",x"99"),
   584 => (x"c0",x"1e",x"cb",x"87"),
   585 => (x"73",x"1e",x"66",x"e0"),
   586 => (x"87",x"e3",x"f1",x"49"),
   587 => (x"98",x"70",x"86",x"c8"),
   588 => (x"87",x"fb",x"c0",x"05"),
   589 => (x"c4",x"4a",x"a3",x"dc"),
   590 => (x"79",x"6a",x"49",x"a4"),
   591 => (x"c8",x"49",x"a3",x"da"),
   592 => (x"69",x"9f",x"4d",x"a4"),
   593 => (x"e0",x"c2",x"7d",x"48"),
   594 => (x"d3",x"02",x"bf",x"c8"),
   595 => (x"49",x"a3",x"d4",x"87"),
   596 => (x"c0",x"49",x"69",x"9f"),
   597 => (x"71",x"99",x"ff",x"ff"),
   598 => (x"c4",x"30",x"d0",x"48"),
   599 => (x"87",x"c2",x"58",x"a6"),
   600 => (x"48",x"6e",x"7e",x"c0"),
   601 => (x"7d",x"70",x"80",x"6d"),
   602 => (x"48",x"c1",x"7c",x"c0"),
   603 => (x"c8",x"87",x"c5",x"c1"),
   604 => (x"80",x"c1",x"48",x"66"),
   605 => (x"c2",x"58",x"a6",x"cc"),
   606 => (x"a8",x"bf",x"cc",x"e0"),
   607 => (x"87",x"e3",x"fd",x"04"),
   608 => (x"bf",x"c8",x"e0",x"c2"),
   609 => (x"87",x"ea",x"c0",x"02"),
   610 => (x"c4",x"fb",x"49",x"6e"),
   611 => (x"58",x"a6",x"c4",x"87"),
   612 => (x"ff",x"cf",x"49",x"70"),
   613 => (x"99",x"f8",x"ff",x"ff"),
   614 => (x"87",x"d6",x"02",x"a9"),
   615 => (x"89",x"c2",x"49",x"70"),
   616 => (x"bf",x"c0",x"e0",x"c2"),
   617 => (x"e0",x"e4",x"c2",x"91"),
   618 => (x"80",x"71",x"48",x"bf"),
   619 => (x"fc",x"58",x"a6",x"c8"),
   620 => (x"48",x"c0",x"87",x"e1"),
   621 => (x"d0",x"f0",x"8e",x"f4"),
   622 => (x"1e",x"73",x"1e",x"87"),
   623 => (x"49",x"6a",x"4a",x"71"),
   624 => (x"7a",x"71",x"81",x"c1"),
   625 => (x"bf",x"c4",x"e0",x"c2"),
   626 => (x"87",x"cb",x"05",x"99"),
   627 => (x"6b",x"4b",x"a2",x"c8"),
   628 => (x"87",x"fd",x"f9",x"49"),
   629 => (x"c1",x"7b",x"49",x"70"),
   630 => (x"87",x"f1",x"ef",x"48"),
   631 => (x"71",x"1e",x"73",x"1e"),
   632 => (x"e0",x"e4",x"c2",x"4b"),
   633 => (x"a3",x"c8",x"49",x"bf"),
   634 => (x"c2",x"4a",x"6a",x"4a"),
   635 => (x"c0",x"e0",x"c2",x"8a"),
   636 => (x"a1",x"72",x"92",x"bf"),
   637 => (x"c4",x"e0",x"c2",x"49"),
   638 => (x"9a",x"6b",x"4a",x"bf"),
   639 => (x"c8",x"49",x"a1",x"72"),
   640 => (x"e8",x"71",x"1e",x"66"),
   641 => (x"86",x"c4",x"87",x"fd"),
   642 => (x"c4",x"05",x"98",x"70"),
   643 => (x"c2",x"48",x"c0",x"87"),
   644 => (x"ee",x"48",x"c1",x"87"),
   645 => (x"5e",x"0e",x"87",x"f7"),
   646 => (x"71",x"0e",x"5c",x"5b"),
   647 => (x"72",x"4b",x"c0",x"4a"),
   648 => (x"e0",x"c0",x"02",x"9a"),
   649 => (x"49",x"a2",x"da",x"87"),
   650 => (x"c2",x"4b",x"69",x"9f"),
   651 => (x"02",x"bf",x"c8",x"e0"),
   652 => (x"a2",x"d4",x"87",x"cf"),
   653 => (x"49",x"69",x"9f",x"49"),
   654 => (x"ff",x"ff",x"c0",x"4c"),
   655 => (x"c2",x"34",x"d0",x"9c"),
   656 => (x"74",x"4c",x"c0",x"87"),
   657 => (x"02",x"9b",x"73",x"b3"),
   658 => (x"c2",x"4a",x"87",x"df"),
   659 => (x"c0",x"e0",x"c2",x"8a"),
   660 => (x"c2",x"92",x"49",x"bf"),
   661 => (x"48",x"bf",x"e0",x"e4"),
   662 => (x"e5",x"c2",x"80",x"72"),
   663 => (x"48",x"71",x"58",x"c0"),
   664 => (x"e0",x"c2",x"30",x"c4"),
   665 => (x"e9",x"c0",x"58",x"d0"),
   666 => (x"e4",x"e4",x"c2",x"87"),
   667 => (x"e4",x"c2",x"4b",x"bf"),
   668 => (x"e4",x"c2",x"48",x"fc"),
   669 => (x"c2",x"78",x"bf",x"e8"),
   670 => (x"02",x"bf",x"c8",x"e0"),
   671 => (x"e0",x"c2",x"87",x"c9"),
   672 => (x"c4",x"49",x"bf",x"c0"),
   673 => (x"c2",x"87",x"c7",x"31"),
   674 => (x"49",x"bf",x"ec",x"e4"),
   675 => (x"e0",x"c2",x"31",x"c4"),
   676 => (x"e4",x"c2",x"59",x"d0"),
   677 => (x"f2",x"ec",x"5b",x"fc"),
   678 => (x"5b",x"5e",x"0e",x"87"),
   679 => (x"f4",x"0e",x"5d",x"5c"),
   680 => (x"9a",x"4a",x"71",x"86"),
   681 => (x"c2",x"87",x"de",x"02"),
   682 => (x"c0",x"48",x"fc",x"d7"),
   683 => (x"f4",x"d7",x"c2",x"78"),
   684 => (x"fc",x"e4",x"c2",x"48"),
   685 => (x"d7",x"c2",x"78",x"bf"),
   686 => (x"e4",x"c2",x"48",x"f8"),
   687 => (x"c0",x"78",x"bf",x"f8"),
   688 => (x"c0",x"48",x"ef",x"f1"),
   689 => (x"cc",x"e0",x"c2",x"78"),
   690 => (x"d7",x"c2",x"49",x"bf"),
   691 => (x"71",x"4a",x"bf",x"fc"),
   692 => (x"cb",x"c4",x"03",x"aa"),
   693 => (x"cf",x"49",x"72",x"87"),
   694 => (x"e0",x"c0",x"05",x"99"),
   695 => (x"c0",x"d8",x"c2",x"87"),
   696 => (x"f4",x"d7",x"c2",x"1e"),
   697 => (x"d7",x"c2",x"49",x"bf"),
   698 => (x"a1",x"c1",x"48",x"f4"),
   699 => (x"d2",x"e5",x"71",x"78"),
   700 => (x"c0",x"86",x"c4",x"87"),
   701 => (x"c2",x"48",x"eb",x"f1"),
   702 => (x"cc",x"78",x"c0",x"d8"),
   703 => (x"eb",x"f1",x"c0",x"87"),
   704 => (x"e0",x"c0",x"48",x"bf"),
   705 => (x"ef",x"f1",x"c0",x"80"),
   706 => (x"fc",x"d7",x"c2",x"58"),
   707 => (x"80",x"c1",x"48",x"bf"),
   708 => (x"58",x"c0",x"d8",x"c2"),
   709 => (x"00",x"0c",x"6b",x"27"),
   710 => (x"bf",x"97",x"bf",x"00"),
   711 => (x"c2",x"02",x"9c",x"4c"),
   712 => (x"e5",x"c3",x"87",x"ee"),
   713 => (x"e7",x"c2",x"02",x"ac"),
   714 => (x"eb",x"f1",x"c0",x"87"),
   715 => (x"a3",x"cb",x"4b",x"bf"),
   716 => (x"cf",x"4d",x"11",x"49"),
   717 => (x"d6",x"c1",x"05",x"ad"),
   718 => (x"df",x"49",x"74",x"87"),
   719 => (x"cd",x"89",x"c1",x"99"),
   720 => (x"d0",x"e0",x"c2",x"91"),
   721 => (x"4a",x"a3",x"c1",x"81"),
   722 => (x"a3",x"c3",x"51",x"12"),
   723 => (x"c5",x"51",x"12",x"4a"),
   724 => (x"51",x"12",x"4a",x"a3"),
   725 => (x"12",x"4a",x"a3",x"c7"),
   726 => (x"4a",x"a3",x"c9",x"51"),
   727 => (x"a3",x"ce",x"51",x"12"),
   728 => (x"d0",x"51",x"12",x"4a"),
   729 => (x"51",x"12",x"4a",x"a3"),
   730 => (x"12",x"4a",x"a3",x"d2"),
   731 => (x"4a",x"a3",x"d4",x"51"),
   732 => (x"a3",x"d6",x"51",x"12"),
   733 => (x"d8",x"51",x"12",x"4a"),
   734 => (x"51",x"12",x"4a",x"a3"),
   735 => (x"12",x"4a",x"a3",x"dc"),
   736 => (x"4a",x"a3",x"de",x"51"),
   737 => (x"f1",x"c0",x"51",x"12"),
   738 => (x"78",x"c1",x"48",x"ef"),
   739 => (x"75",x"87",x"c1",x"c1"),
   740 => (x"05",x"99",x"c8",x"49"),
   741 => (x"75",x"87",x"f3",x"c0"),
   742 => (x"05",x"99",x"d0",x"49"),
   743 => (x"66",x"dc",x"87",x"d0"),
   744 => (x"87",x"ca",x"c0",x"02"),
   745 => (x"66",x"dc",x"49",x"73"),
   746 => (x"02",x"98",x"70",x"0f"),
   747 => (x"f1",x"c0",x"87",x"dc"),
   748 => (x"c0",x"05",x"bf",x"ef"),
   749 => (x"e0",x"c2",x"87",x"c6"),
   750 => (x"50",x"c0",x"48",x"d0"),
   751 => (x"48",x"ef",x"f1",x"c0"),
   752 => (x"f1",x"c0",x"78",x"c0"),
   753 => (x"c2",x"48",x"bf",x"eb"),
   754 => (x"f1",x"c0",x"87",x"dc"),
   755 => (x"78",x"c0",x"48",x"ef"),
   756 => (x"bf",x"cc",x"e0",x"c2"),
   757 => (x"fc",x"d7",x"c2",x"49"),
   758 => (x"aa",x"71",x"4a",x"bf"),
   759 => (x"87",x"f5",x"fb",x"04"),
   760 => (x"bf",x"fc",x"e4",x"c2"),
   761 => (x"87",x"c8",x"c0",x"05"),
   762 => (x"bf",x"c8",x"e0",x"c2"),
   763 => (x"87",x"f4",x"c1",x"02"),
   764 => (x"bf",x"f8",x"d7",x"c2"),
   765 => (x"87",x"d9",x"f1",x"49"),
   766 => (x"58",x"fc",x"d7",x"c2"),
   767 => (x"e0",x"c2",x"7e",x"70"),
   768 => (x"c0",x"02",x"bf",x"c8"),
   769 => (x"49",x"6e",x"87",x"dd"),
   770 => (x"ff",x"ff",x"ff",x"cf"),
   771 => (x"02",x"a9",x"99",x"f8"),
   772 => (x"c4",x"87",x"c8",x"c0"),
   773 => (x"78",x"c0",x"48",x"a6"),
   774 => (x"c4",x"87",x"e6",x"c0"),
   775 => (x"78",x"c1",x"48",x"a6"),
   776 => (x"6e",x"87",x"de",x"c0"),
   777 => (x"f8",x"ff",x"cf",x"49"),
   778 => (x"c0",x"02",x"a9",x"99"),
   779 => (x"a6",x"c8",x"87",x"c8"),
   780 => (x"c0",x"78",x"c0",x"48"),
   781 => (x"a6",x"c8",x"87",x"c5"),
   782 => (x"c4",x"78",x"c1",x"48"),
   783 => (x"66",x"c8",x"48",x"a6"),
   784 => (x"05",x"66",x"c4",x"78"),
   785 => (x"6e",x"87",x"dd",x"c0"),
   786 => (x"c2",x"89",x"c2",x"49"),
   787 => (x"91",x"bf",x"c0",x"e0"),
   788 => (x"bf",x"e0",x"e4",x"c2"),
   789 => (x"c2",x"80",x"71",x"48"),
   790 => (x"c2",x"58",x"f8",x"d7"),
   791 => (x"c0",x"48",x"fc",x"d7"),
   792 => (x"87",x"e1",x"f9",x"78"),
   793 => (x"8e",x"f4",x"48",x"c0"),
   794 => (x"00",x"87",x"de",x"e5"),
   795 => (x"00",x"00",x"00",x"00"),
   796 => (x"1e",x"00",x"00",x"00"),
   797 => (x"c3",x"48",x"d4",x"ff"),
   798 => (x"49",x"68",x"78",x"ff"),
   799 => (x"87",x"c6",x"02",x"99"),
   800 => (x"05",x"a9",x"fb",x"c0"),
   801 => (x"48",x"71",x"87",x"ee"),
   802 => (x"5e",x"0e",x"4f",x"26"),
   803 => (x"71",x"0e",x"5c",x"5b"),
   804 => (x"ff",x"4b",x"c0",x"4a"),
   805 => (x"ff",x"c3",x"48",x"d4"),
   806 => (x"99",x"49",x"68",x"78"),
   807 => (x"87",x"c1",x"c1",x"02"),
   808 => (x"02",x"a9",x"ec",x"c0"),
   809 => (x"c0",x"87",x"fa",x"c0"),
   810 => (x"c0",x"02",x"a9",x"fb"),
   811 => (x"66",x"cc",x"87",x"f3"),
   812 => (x"cc",x"03",x"ab",x"b7"),
   813 => (x"02",x"66",x"d0",x"87"),
   814 => (x"09",x"72",x"87",x"c7"),
   815 => (x"c1",x"09",x"79",x"97"),
   816 => (x"02",x"99",x"71",x"82"),
   817 => (x"83",x"c1",x"87",x"c2"),
   818 => (x"c3",x"48",x"d4",x"ff"),
   819 => (x"49",x"68",x"78",x"ff"),
   820 => (x"87",x"cd",x"02",x"99"),
   821 => (x"02",x"a9",x"ec",x"c0"),
   822 => (x"fb",x"c0",x"87",x"c7"),
   823 => (x"cd",x"ff",x"05",x"a9"),
   824 => (x"02",x"66",x"d0",x"87"),
   825 => (x"97",x"c0",x"87",x"c3"),
   826 => (x"a9",x"fb",x"c0",x"7a"),
   827 => (x"73",x"87",x"c7",x"05"),
   828 => (x"8c",x"0c",x"c0",x"4c"),
   829 => (x"4c",x"73",x"87",x"c2"),
   830 => (x"87",x"c2",x"48",x"74"),
   831 => (x"4c",x"26",x"4d",x"26"),
   832 => (x"4f",x"26",x"4b",x"26"),
   833 => (x"48",x"d4",x"ff",x"1e"),
   834 => (x"68",x"78",x"ff",x"c3"),
   835 => (x"b7",x"f0",x"c0",x"49"),
   836 => (x"87",x"ca",x"04",x"a9"),
   837 => (x"a9",x"b7",x"f9",x"c0"),
   838 => (x"c0",x"87",x"c3",x"01"),
   839 => (x"c1",x"c1",x"89",x"f0"),
   840 => (x"ca",x"04",x"a9",x"b7"),
   841 => (x"b7",x"c6",x"c1",x"87"),
   842 => (x"87",x"c3",x"01",x"a9"),
   843 => (x"71",x"89",x"f7",x"c0"),
   844 => (x"0e",x"4f",x"26",x"48"),
   845 => (x"5d",x"5c",x"5b",x"5e"),
   846 => (x"71",x"86",x"f4",x"0e"),
   847 => (x"4b",x"d4",x"ff",x"4c"),
   848 => (x"c3",x"7e",x"4d",x"c0"),
   849 => (x"d0",x"ff",x"7b",x"ff"),
   850 => (x"c0",x"c8",x"48",x"bf"),
   851 => (x"a6",x"c8",x"98",x"c0"),
   852 => (x"02",x"98",x"70",x"58"),
   853 => (x"d0",x"ff",x"87",x"d0"),
   854 => (x"c0",x"c8",x"48",x"bf"),
   855 => (x"a6",x"c8",x"98",x"c0"),
   856 => (x"05",x"98",x"70",x"58"),
   857 => (x"d0",x"ff",x"87",x"f0"),
   858 => (x"78",x"e1",x"c0",x"48"),
   859 => (x"c2",x"fc",x"7b",x"d4"),
   860 => (x"99",x"49",x"70",x"87"),
   861 => (x"87",x"c7",x"c1",x"02"),
   862 => (x"c8",x"7b",x"ff",x"c3"),
   863 => (x"78",x"6b",x"48",x"a6"),
   864 => (x"c0",x"48",x"66",x"c8"),
   865 => (x"c8",x"02",x"a8",x"fb"),
   866 => (x"d8",x"e5",x"c2",x"87"),
   867 => (x"ee",x"c0",x"02",x"bf"),
   868 => (x"71",x"4d",x"c1",x"87"),
   869 => (x"e6",x"c0",x"02",x"99"),
   870 => (x"a9",x"fb",x"c0",x"87"),
   871 => (x"fb",x"87",x"c3",x"02"),
   872 => (x"ff",x"c3",x"87",x"d1"),
   873 => (x"c1",x"49",x"6b",x"7b"),
   874 => (x"cc",x"05",x"a9",x"c6"),
   875 => (x"7b",x"ff",x"c3",x"87"),
   876 => (x"48",x"a6",x"c8",x"7b"),
   877 => (x"49",x"c0",x"78",x"6b"),
   878 => (x"05",x"99",x"71",x"4d"),
   879 => (x"75",x"87",x"da",x"ff"),
   880 => (x"de",x"c1",x"05",x"9d"),
   881 => (x"7b",x"ff",x"c3",x"87"),
   882 => (x"ff",x"c3",x"4a",x"6b"),
   883 => (x"48",x"a6",x"c4",x"7b"),
   884 => (x"48",x"6e",x"78",x"6b"),
   885 => (x"a6",x"c4",x"80",x"c1"),
   886 => (x"49",x"a4",x"c8",x"58"),
   887 => (x"c8",x"49",x"69",x"97"),
   888 => (x"da",x"05",x"a9",x"66"),
   889 => (x"49",x"a4",x"c9",x"87"),
   890 => (x"aa",x"49",x"69",x"97"),
   891 => (x"ca",x"87",x"d0",x"05"),
   892 => (x"69",x"97",x"49",x"a4"),
   893 => (x"a9",x"66",x"c4",x"49"),
   894 => (x"c1",x"87",x"c4",x"05"),
   895 => (x"c8",x"87",x"d6",x"4d"),
   896 => (x"ec",x"c0",x"48",x"66"),
   897 => (x"87",x"c9",x"02",x"a8"),
   898 => (x"c0",x"48",x"66",x"c8"),
   899 => (x"c4",x"05",x"a8",x"fb"),
   900 => (x"c1",x"7e",x"c0",x"87"),
   901 => (x"7b",x"ff",x"c3",x"4d"),
   902 => (x"6b",x"48",x"a6",x"c8"),
   903 => (x"02",x"9d",x"75",x"78"),
   904 => (x"ff",x"87",x"e2",x"fe"),
   905 => (x"c8",x"48",x"bf",x"d0"),
   906 => (x"c8",x"98",x"c0",x"c0"),
   907 => (x"98",x"70",x"58",x"a6"),
   908 => (x"ff",x"87",x"d0",x"02"),
   909 => (x"c8",x"48",x"bf",x"d0"),
   910 => (x"c8",x"98",x"c0",x"c0"),
   911 => (x"98",x"70",x"58",x"a6"),
   912 => (x"ff",x"87",x"f0",x"05"),
   913 => (x"e0",x"c0",x"48",x"d0"),
   914 => (x"f4",x"48",x"6e",x"78"),
   915 => (x"87",x"ec",x"fa",x"8e"),
   916 => (x"5c",x"5b",x"5e",x"0e"),
   917 => (x"86",x"f4",x"0e",x"5d"),
   918 => (x"ff",x"59",x"a6",x"c4"),
   919 => (x"c0",x"c8",x"4c",x"d0"),
   920 => (x"1e",x"6e",x"4b",x"c0"),
   921 => (x"49",x"dc",x"e5",x"c2"),
   922 => (x"c4",x"87",x"cf",x"e9"),
   923 => (x"02",x"98",x"70",x"86"),
   924 => (x"c2",x"87",x"f7",x"c5"),
   925 => (x"4d",x"bf",x"e0",x"e5"),
   926 => (x"f6",x"fa",x"49",x"6e"),
   927 => (x"58",x"a6",x"c8",x"87"),
   928 => (x"98",x"73",x"48",x"6c"),
   929 => (x"70",x"58",x"a6",x"cc"),
   930 => (x"87",x"cc",x"02",x"98"),
   931 => (x"98",x"73",x"48",x"6c"),
   932 => (x"70",x"58",x"a6",x"c4"),
   933 => (x"87",x"f4",x"05",x"98"),
   934 => (x"d4",x"ff",x"7c",x"c5"),
   935 => (x"78",x"d5",x"c1",x"48"),
   936 => (x"bf",x"d8",x"e5",x"c2"),
   937 => (x"c4",x"81",x"c1",x"49"),
   938 => (x"8a",x"c1",x"4a",x"66"),
   939 => (x"48",x"72",x"32",x"c6"),
   940 => (x"d4",x"ff",x"b0",x"71"),
   941 => (x"48",x"6c",x"78",x"08"),
   942 => (x"a6",x"c4",x"98",x"73"),
   943 => (x"02",x"98",x"70",x"58"),
   944 => (x"48",x"6c",x"87",x"cc"),
   945 => (x"a6",x"c4",x"98",x"73"),
   946 => (x"05",x"98",x"70",x"58"),
   947 => (x"7c",x"c4",x"87",x"f4"),
   948 => (x"c3",x"48",x"d4",x"ff"),
   949 => (x"48",x"6c",x"78",x"ff"),
   950 => (x"a6",x"c4",x"98",x"73"),
   951 => (x"02",x"98",x"70",x"58"),
   952 => (x"48",x"6c",x"87",x"cc"),
   953 => (x"a6",x"c4",x"98",x"73"),
   954 => (x"05",x"98",x"70",x"58"),
   955 => (x"7c",x"c5",x"87",x"f4"),
   956 => (x"c1",x"48",x"d4",x"ff"),
   957 => (x"78",x"c1",x"78",x"d3"),
   958 => (x"98",x"73",x"48",x"6c"),
   959 => (x"70",x"58",x"a6",x"c4"),
   960 => (x"87",x"cc",x"02",x"98"),
   961 => (x"98",x"73",x"48",x"6c"),
   962 => (x"70",x"58",x"a6",x"c4"),
   963 => (x"87",x"f4",x"05",x"98"),
   964 => (x"9d",x"75",x"7c",x"c4"),
   965 => (x"87",x"d0",x"c2",x"02"),
   966 => (x"7e",x"c0",x"d8",x"c2"),
   967 => (x"dc",x"e5",x"c2",x"1e"),
   968 => (x"87",x"f8",x"ea",x"49"),
   969 => (x"98",x"70",x"86",x"c4"),
   970 => (x"c0",x"87",x"c5",x"05"),
   971 => (x"87",x"fc",x"c2",x"48"),
   972 => (x"ad",x"b7",x"c0",x"c8"),
   973 => (x"4a",x"87",x"c4",x"04"),
   974 => (x"75",x"87",x"c4",x"8d"),
   975 => (x"6c",x"4d",x"c0",x"4a"),
   976 => (x"c8",x"98",x"73",x"48"),
   977 => (x"98",x"70",x"58",x"a6"),
   978 => (x"6c",x"87",x"cc",x"02"),
   979 => (x"c8",x"98",x"73",x"48"),
   980 => (x"98",x"70",x"58",x"a6"),
   981 => (x"cd",x"87",x"f4",x"05"),
   982 => (x"48",x"d4",x"ff",x"7c"),
   983 => (x"72",x"78",x"d4",x"c1"),
   984 => (x"71",x"8a",x"c1",x"49"),
   985 => (x"87",x"d9",x"02",x"99"),
   986 => (x"48",x"bf",x"97",x"6e"),
   987 => (x"78",x"08",x"d4",x"ff"),
   988 => (x"80",x"c1",x"48",x"6e"),
   989 => (x"72",x"58",x"a6",x"c4"),
   990 => (x"71",x"8a",x"c1",x"49"),
   991 => (x"e7",x"ff",x"05",x"99"),
   992 => (x"73",x"48",x"6c",x"87"),
   993 => (x"58",x"a6",x"c4",x"98"),
   994 => (x"cc",x"02",x"98",x"70"),
   995 => (x"73",x"48",x"6c",x"87"),
   996 => (x"58",x"a6",x"c4",x"98"),
   997 => (x"f4",x"05",x"98",x"70"),
   998 => (x"c2",x"7c",x"c4",x"87"),
   999 => (x"e8",x"49",x"dc",x"e5"),
  1000 => (x"9d",x"75",x"87",x"d7"),
  1001 => (x"87",x"f0",x"fd",x"05"),
  1002 => (x"98",x"73",x"48",x"6c"),
  1003 => (x"70",x"58",x"a6",x"c4"),
  1004 => (x"87",x"cd",x"02",x"98"),
  1005 => (x"98",x"73",x"48",x"6c"),
  1006 => (x"70",x"58",x"a6",x"c4"),
  1007 => (x"f3",x"ff",x"05",x"98"),
  1008 => (x"ff",x"7c",x"c5",x"87"),
  1009 => (x"d3",x"c1",x"48",x"d4"),
  1010 => (x"6c",x"78",x"c0",x"78"),
  1011 => (x"c4",x"98",x"73",x"48"),
  1012 => (x"98",x"70",x"58",x"a6"),
  1013 => (x"6c",x"87",x"cd",x"02"),
  1014 => (x"c4",x"98",x"73",x"48"),
  1015 => (x"98",x"70",x"58",x"a6"),
  1016 => (x"87",x"f3",x"ff",x"05"),
  1017 => (x"48",x"c1",x"7c",x"c4"),
  1018 => (x"48",x"c0",x"87",x"c2"),
  1019 => (x"cb",x"f4",x"8e",x"f4"),
  1020 => (x"5b",x"5e",x"0e",x"87"),
  1021 => (x"1e",x"0e",x"5d",x"5c"),
  1022 => (x"4c",x"c0",x"4b",x"71"),
  1023 => (x"04",x"ab",x"b7",x"4d"),
  1024 => (x"c0",x"87",x"e9",x"c0"),
  1025 => (x"75",x"1e",x"f3",x"f4"),
  1026 => (x"87",x"c4",x"02",x"9d"),
  1027 => (x"87",x"c2",x"4a",x"c0"),
  1028 => (x"49",x"72",x"4a",x"c1"),
  1029 => (x"c4",x"87",x"c2",x"ea"),
  1030 => (x"c1",x"58",x"a6",x"86"),
  1031 => (x"c2",x"05",x"6e",x"84"),
  1032 => (x"c1",x"4c",x"73",x"87"),
  1033 => (x"ac",x"b7",x"73",x"85"),
  1034 => (x"87",x"d7",x"ff",x"06"),
  1035 => (x"f3",x"26",x"48",x"6e"),
  1036 => (x"5e",x"0e",x"87",x"ca"),
  1037 => (x"0e",x"5d",x"5c",x"5b"),
  1038 => (x"49",x"4c",x"71",x"1e"),
  1039 => (x"bf",x"ec",x"e5",x"c2"),
  1040 => (x"87",x"ed",x"fe",x"81"),
  1041 => (x"02",x"9d",x"4d",x"70"),
  1042 => (x"c2",x"87",x"fc",x"c0"),
  1043 => (x"75",x"4b",x"d0",x"e0"),
  1044 => (x"ff",x"49",x"cb",x"4a"),
  1045 => (x"74",x"87",x"c9",x"c1"),
  1046 => (x"c2",x"91",x"de",x"49"),
  1047 => (x"71",x"48",x"c0",x"e6"),
  1048 => (x"58",x"a6",x"c4",x"80"),
  1049 => (x"48",x"d7",x"c2",x"c1"),
  1050 => (x"a1",x"c8",x"49",x"6e"),
  1051 => (x"71",x"41",x"20",x"4a"),
  1052 => (x"87",x"f9",x"05",x"aa"),
  1053 => (x"51",x"10",x"51",x"10"),
  1054 => (x"49",x"74",x"51",x"10"),
  1055 => (x"87",x"ee",x"c5",x"c1"),
  1056 => (x"49",x"d0",x"e0",x"c2"),
  1057 => (x"c1",x"87",x"c9",x"f7"),
  1058 => (x"c1",x"49",x"d0",x"e4"),
  1059 => (x"c1",x"87",x"f6",x"c7"),
  1060 => (x"26",x"87",x"d2",x"c8"),
  1061 => (x"4c",x"87",x"e5",x"f1"),
  1062 => (x"69",x"64",x"61",x"6f"),
  1063 => (x"2e",x"2e",x"67",x"6e"),
  1064 => (x"20",x"80",x"00",x"2e"),
  1065 => (x"6b",x"63",x"61",x"42"),
  1066 => (x"61",x"6f",x"4c",x"00"),
  1067 => (x"2e",x"2a",x"20",x"64"),
  1068 => (x"20",x"3a",x"00",x"20"),
  1069 => (x"42",x"20",x"80",x"00"),
  1070 => (x"00",x"6b",x"63",x"61"),
  1071 => (x"78",x"45",x"20",x"80"),
  1072 => (x"53",x"00",x"74",x"69"),
  1073 => (x"6e",x"49",x"20",x"44"),
  1074 => (x"2e",x"2e",x"74",x"69"),
  1075 => (x"00",x"4b",x"4f",x"00"),
  1076 => (x"54",x"4f",x"4f",x"42"),
  1077 => (x"20",x"20",x"20",x"20"),
  1078 => (x"00",x"4d",x"4f",x"52"),
  1079 => (x"71",x"1e",x"73",x"1e"),
  1080 => (x"e5",x"c2",x"49",x"4b"),
  1081 => (x"fc",x"81",x"bf",x"ec"),
  1082 => (x"4a",x"70",x"87",x"c7"),
  1083 => (x"87",x"c4",x"02",x"9a"),
  1084 => (x"87",x"e2",x"e4",x"49"),
  1085 => (x"48",x"ec",x"e5",x"c2"),
  1086 => (x"49",x"73",x"78",x"c0"),
  1087 => (x"ef",x"87",x"e9",x"c1"),
  1088 => (x"73",x"1e",x"87",x"fe"),
  1089 => (x"c4",x"4b",x"71",x"1e"),
  1090 => (x"c1",x"02",x"4a",x"a3"),
  1091 => (x"8a",x"c1",x"87",x"c8"),
  1092 => (x"8a",x"87",x"dc",x"02"),
  1093 => (x"87",x"f1",x"c0",x"02"),
  1094 => (x"c4",x"c1",x"05",x"8a"),
  1095 => (x"ec",x"e5",x"c2",x"87"),
  1096 => (x"fc",x"c0",x"02",x"bf"),
  1097 => (x"88",x"c1",x"48",x"87"),
  1098 => (x"58",x"f0",x"e5",x"c2"),
  1099 => (x"c2",x"87",x"f2",x"c0"),
  1100 => (x"49",x"bf",x"ec",x"e5"),
  1101 => (x"e5",x"c2",x"89",x"d0"),
  1102 => (x"b7",x"c0",x"59",x"f0"),
  1103 => (x"e0",x"c0",x"03",x"a9"),
  1104 => (x"ec",x"e5",x"c2",x"87"),
  1105 => (x"d8",x"78",x"c0",x"48"),
  1106 => (x"ec",x"e5",x"c2",x"87"),
  1107 => (x"80",x"c1",x"48",x"bf"),
  1108 => (x"58",x"f0",x"e5",x"c2"),
  1109 => (x"e5",x"c2",x"87",x"cb"),
  1110 => (x"d0",x"48",x"bf",x"ec"),
  1111 => (x"f0",x"e5",x"c2",x"80"),
  1112 => (x"c3",x"49",x"73",x"58"),
  1113 => (x"87",x"d8",x"ee",x"87"),
  1114 => (x"5c",x"5b",x"5e",x"0e"),
  1115 => (x"86",x"f0",x"0e",x"5d"),
  1116 => (x"c2",x"59",x"a6",x"d0"),
  1117 => (x"c0",x"4d",x"c0",x"d8"),
  1118 => (x"48",x"a6",x"c4",x"4c"),
  1119 => (x"e5",x"c2",x"78",x"c0"),
  1120 => (x"c0",x"48",x"bf",x"ec"),
  1121 => (x"c1",x"06",x"a8",x"b7"),
  1122 => (x"d8",x"c2",x"87",x"c1"),
  1123 => (x"02",x"98",x"48",x"c0"),
  1124 => (x"c0",x"87",x"f8",x"c0"),
  1125 => (x"c8",x"1e",x"f3",x"f4"),
  1126 => (x"87",x"c7",x"02",x"66"),
  1127 => (x"c0",x"48",x"a6",x"c4"),
  1128 => (x"c4",x"87",x"c5",x"78"),
  1129 => (x"78",x"c1",x"48",x"a6"),
  1130 => (x"e3",x"49",x"66",x"c4"),
  1131 => (x"86",x"c4",x"87",x"eb"),
  1132 => (x"84",x"c1",x"4d",x"70"),
  1133 => (x"c1",x"48",x"66",x"c4"),
  1134 => (x"58",x"a6",x"c8",x"80"),
  1135 => (x"bf",x"ec",x"e5",x"c2"),
  1136 => (x"c6",x"03",x"ac",x"b7"),
  1137 => (x"05",x"9d",x"75",x"87"),
  1138 => (x"c0",x"87",x"c8",x"ff"),
  1139 => (x"02",x"9d",x"75",x"4c"),
  1140 => (x"c0",x"87",x"e3",x"c3"),
  1141 => (x"c8",x"1e",x"f3",x"f4"),
  1142 => (x"87",x"c7",x"02",x"66"),
  1143 => (x"c0",x"48",x"a6",x"cc"),
  1144 => (x"cc",x"87",x"c5",x"78"),
  1145 => (x"78",x"c1",x"48",x"a6"),
  1146 => (x"e2",x"49",x"66",x"cc"),
  1147 => (x"86",x"c4",x"87",x"eb"),
  1148 => (x"02",x"6e",x"58",x"a6"),
  1149 => (x"49",x"87",x"eb",x"c2"),
  1150 => (x"69",x"97",x"81",x"cb"),
  1151 => (x"02",x"99",x"d0",x"49"),
  1152 => (x"c1",x"87",x"d9",x"c1"),
  1153 => (x"74",x"4b",x"dc",x"c3"),
  1154 => (x"c1",x"91",x"cc",x"49"),
  1155 => (x"c8",x"81",x"d0",x"e4"),
  1156 => (x"7a",x"73",x"4a",x"a1"),
  1157 => (x"ff",x"c3",x"81",x"c1"),
  1158 => (x"de",x"49",x"74",x"51"),
  1159 => (x"c0",x"e6",x"c2",x"91"),
  1160 => (x"c2",x"85",x"71",x"4d"),
  1161 => (x"c1",x"7d",x"97",x"c1"),
  1162 => (x"e0",x"c0",x"49",x"a5"),
  1163 => (x"d0",x"e0",x"c2",x"51"),
  1164 => (x"d2",x"02",x"bf",x"97"),
  1165 => (x"c2",x"84",x"c1",x"87"),
  1166 => (x"e0",x"c2",x"4b",x"a5"),
  1167 => (x"49",x"db",x"4a",x"d0"),
  1168 => (x"87",x"dc",x"f9",x"fe"),
  1169 => (x"cd",x"87",x"db",x"c1"),
  1170 => (x"51",x"c0",x"49",x"a5"),
  1171 => (x"a5",x"c2",x"84",x"c1"),
  1172 => (x"cb",x"4a",x"6e",x"4b"),
  1173 => (x"c7",x"f9",x"fe",x"49"),
  1174 => (x"87",x"c6",x"c1",x"87"),
  1175 => (x"91",x"cc",x"49",x"74"),
  1176 => (x"81",x"d0",x"e4",x"c1"),
  1177 => (x"c0",x"c1",x"81",x"c8"),
  1178 => (x"e0",x"c2",x"79",x"f2"),
  1179 => (x"02",x"bf",x"97",x"d0"),
  1180 => (x"49",x"74",x"87",x"d8"),
  1181 => (x"84",x"c1",x"91",x"de"),
  1182 => (x"4b",x"c0",x"e6",x"c2"),
  1183 => (x"e0",x"c2",x"83",x"71"),
  1184 => (x"49",x"dd",x"4a",x"d0"),
  1185 => (x"87",x"d8",x"f8",x"fe"),
  1186 => (x"4b",x"74",x"87",x"d8"),
  1187 => (x"e6",x"c2",x"93",x"de"),
  1188 => (x"a3",x"cb",x"83",x"c0"),
  1189 => (x"c1",x"51",x"c0",x"49"),
  1190 => (x"4a",x"6e",x"73",x"84"),
  1191 => (x"f7",x"fe",x"49",x"cb"),
  1192 => (x"66",x"c4",x"87",x"fe"),
  1193 => (x"c8",x"80",x"c1",x"48"),
  1194 => (x"b7",x"c7",x"58",x"a6"),
  1195 => (x"c5",x"c0",x"03",x"ac"),
  1196 => (x"fc",x"05",x"6e",x"87"),
  1197 => (x"b7",x"c7",x"87",x"dd"),
  1198 => (x"d3",x"c0",x"03",x"ac"),
  1199 => (x"de",x"49",x"74",x"87"),
  1200 => (x"c0",x"e6",x"c2",x"91"),
  1201 => (x"c1",x"51",x"c0",x"81"),
  1202 => (x"ac",x"b7",x"c7",x"84"),
  1203 => (x"87",x"ed",x"ff",x"04"),
  1204 => (x"48",x"e5",x"e5",x"c1"),
  1205 => (x"e5",x"c1",x"50",x"c0"),
  1206 => (x"50",x"c2",x"48",x"e4"),
  1207 => (x"48",x"ec",x"e5",x"c1"),
  1208 => (x"78",x"ce",x"cc",x"c1"),
  1209 => (x"48",x"e8",x"e5",x"c1"),
  1210 => (x"78",x"e2",x"c2",x"c1"),
  1211 => (x"48",x"f8",x"e5",x"c1"),
  1212 => (x"78",x"c2",x"c4",x"c1"),
  1213 => (x"c0",x"49",x"66",x"cc"),
  1214 => (x"f0",x"87",x"f3",x"fb"),
  1215 => (x"87",x"fc",x"e7",x"8e"),
  1216 => (x"c2",x"4a",x"71",x"1e"),
  1217 => (x"72",x"5a",x"dc",x"e5"),
  1218 => (x"87",x"dc",x"f9",x"49"),
  1219 => (x"71",x"1e",x"4f",x"26"),
  1220 => (x"91",x"cc",x"49",x"4a"),
  1221 => (x"81",x"d0",x"e4",x"c1"),
  1222 => (x"48",x"11",x"81",x"c1"),
  1223 => (x"58",x"d8",x"e5",x"c2"),
  1224 => (x"49",x"a2",x"f0",x"c0"),
  1225 => (x"87",x"c8",x"f6",x"fe"),
  1226 => (x"dd",x"d5",x"49",x"c0"),
  1227 => (x"0e",x"4f",x"26",x"87"),
  1228 => (x"5d",x"5c",x"5b",x"5e"),
  1229 => (x"71",x"86",x"f0",x"0e"),
  1230 => (x"91",x"cc",x"49",x"4c"),
  1231 => (x"81",x"d0",x"e4",x"c1"),
  1232 => (x"c4",x"7e",x"a1",x"c3"),
  1233 => (x"e5",x"c2",x"48",x"a6"),
  1234 => (x"6e",x"78",x"bf",x"d0"),
  1235 => (x"c4",x"4a",x"bf",x"97"),
  1236 => (x"2b",x"72",x"4b",x"66"),
  1237 => (x"12",x"4a",x"a1",x"c1"),
  1238 => (x"58",x"a6",x"cc",x"48"),
  1239 => (x"83",x"c1",x"9b",x"70"),
  1240 => (x"69",x"97",x"81",x"c2"),
  1241 => (x"04",x"ab",x"b7",x"49"),
  1242 => (x"4b",x"c0",x"87",x"c2"),
  1243 => (x"4a",x"bf",x"97",x"6e"),
  1244 => (x"72",x"49",x"66",x"c8"),
  1245 => (x"c4",x"b9",x"ff",x"31"),
  1246 => (x"4d",x"73",x"99",x"66"),
  1247 => (x"b5",x"71",x"35",x"72"),
  1248 => (x"5d",x"d4",x"e5",x"c2"),
  1249 => (x"c3",x"48",x"d4",x"ff"),
  1250 => (x"d0",x"ff",x"78",x"ff"),
  1251 => (x"c0",x"c8",x"48",x"bf"),
  1252 => (x"a6",x"d0",x"98",x"c0"),
  1253 => (x"02",x"98",x"70",x"58"),
  1254 => (x"d0",x"ff",x"87",x"d0"),
  1255 => (x"c0",x"c8",x"48",x"bf"),
  1256 => (x"a6",x"c4",x"98",x"c0"),
  1257 => (x"05",x"98",x"70",x"58"),
  1258 => (x"d0",x"ff",x"87",x"f0"),
  1259 => (x"78",x"e1",x"c0",x"48"),
  1260 => (x"de",x"48",x"d4",x"ff"),
  1261 => (x"7d",x"0d",x"70",x"78"),
  1262 => (x"c8",x"48",x"75",x"0d"),
  1263 => (x"d4",x"ff",x"28",x"b7"),
  1264 => (x"48",x"75",x"78",x"08"),
  1265 => (x"ff",x"28",x"b7",x"d0"),
  1266 => (x"75",x"78",x"08",x"d4"),
  1267 => (x"28",x"b7",x"d8",x"48"),
  1268 => (x"78",x"08",x"d4",x"ff"),
  1269 => (x"48",x"bf",x"d0",x"ff"),
  1270 => (x"98",x"c0",x"c0",x"c8"),
  1271 => (x"70",x"58",x"a6",x"c4"),
  1272 => (x"87",x"d0",x"02",x"98"),
  1273 => (x"48",x"bf",x"d0",x"ff"),
  1274 => (x"98",x"c0",x"c0",x"c8"),
  1275 => (x"70",x"58",x"a6",x"c4"),
  1276 => (x"87",x"f0",x"05",x"98"),
  1277 => (x"c0",x"48",x"d0",x"ff"),
  1278 => (x"1e",x"c7",x"78",x"e0"),
  1279 => (x"e4",x"c1",x"1e",x"c0"),
  1280 => (x"e5",x"c2",x"1e",x"d0"),
  1281 => (x"c1",x"49",x"bf",x"d4"),
  1282 => (x"49",x"74",x"87",x"e1"),
  1283 => (x"87",x"de",x"f7",x"c0"),
  1284 => (x"e7",x"e3",x"8e",x"e4"),
  1285 => (x"1e",x"73",x"1e",x"87"),
  1286 => (x"fc",x"49",x"4b",x"71"),
  1287 => (x"49",x"73",x"87",x"d1"),
  1288 => (x"e3",x"87",x"cc",x"fc"),
  1289 => (x"73",x"1e",x"87",x"da"),
  1290 => (x"c2",x"4b",x"71",x"1e"),
  1291 => (x"d5",x"02",x"4a",x"a3"),
  1292 => (x"05",x"8a",x"c1",x"87"),
  1293 => (x"e5",x"c2",x"87",x"db"),
  1294 => (x"d4",x"02",x"bf",x"e8"),
  1295 => (x"88",x"c1",x"48",x"87"),
  1296 => (x"58",x"ec",x"e5",x"c2"),
  1297 => (x"e5",x"c2",x"87",x"cb"),
  1298 => (x"c1",x"48",x"bf",x"e8"),
  1299 => (x"ec",x"e5",x"c2",x"80"),
  1300 => (x"c0",x"1e",x"c7",x"58"),
  1301 => (x"d0",x"e4",x"c1",x"1e"),
  1302 => (x"d4",x"e5",x"c2",x"1e"),
  1303 => (x"87",x"cb",x"49",x"bf"),
  1304 => (x"f6",x"c0",x"49",x"73"),
  1305 => (x"8e",x"f4",x"87",x"c8"),
  1306 => (x"0e",x"87",x"d5",x"e2"),
  1307 => (x"5d",x"5c",x"5b",x"5e"),
  1308 => (x"86",x"d8",x"ff",x"0e"),
  1309 => (x"c8",x"59",x"a6",x"dc"),
  1310 => (x"78",x"c0",x"48",x"a6"),
  1311 => (x"78",x"c0",x"80",x"c4"),
  1312 => (x"c2",x"80",x"c4",x"4d"),
  1313 => (x"78",x"bf",x"e8",x"e5"),
  1314 => (x"c3",x"48",x"d4",x"ff"),
  1315 => (x"d0",x"ff",x"78",x"ff"),
  1316 => (x"c0",x"c8",x"48",x"bf"),
  1317 => (x"a6",x"c4",x"98",x"c0"),
  1318 => (x"02",x"98",x"70",x"58"),
  1319 => (x"d0",x"ff",x"87",x"d0"),
  1320 => (x"c0",x"c8",x"48",x"bf"),
  1321 => (x"a6",x"c4",x"98",x"c0"),
  1322 => (x"05",x"98",x"70",x"58"),
  1323 => (x"d0",x"ff",x"87",x"f0"),
  1324 => (x"78",x"e1",x"c0",x"48"),
  1325 => (x"d4",x"48",x"d4",x"ff"),
  1326 => (x"f6",x"de",x"ff",x"78"),
  1327 => (x"48",x"d4",x"ff",x"87"),
  1328 => (x"d4",x"78",x"ff",x"c3"),
  1329 => (x"d4",x"ff",x"48",x"a6"),
  1330 => (x"66",x"d4",x"78",x"bf"),
  1331 => (x"a8",x"fb",x"c0",x"48"),
  1332 => (x"87",x"d3",x"c1",x"02"),
  1333 => (x"4a",x"66",x"f8",x"c0"),
  1334 => (x"7e",x"6a",x"82",x"c4"),
  1335 => (x"c2",x"c1",x"1e",x"72"),
  1336 => (x"66",x"c4",x"48",x"e9"),
  1337 => (x"4a",x"a1",x"c8",x"49"),
  1338 => (x"aa",x"71",x"41",x"20"),
  1339 => (x"10",x"87",x"f9",x"05"),
  1340 => (x"c0",x"4a",x"26",x"51"),
  1341 => (x"c8",x"49",x"66",x"f8"),
  1342 => (x"c0",x"cc",x"c1",x"81"),
  1343 => (x"c7",x"49",x"6a",x"79"),
  1344 => (x"51",x"66",x"d4",x"81"),
  1345 => (x"1e",x"d8",x"1e",x"c1"),
  1346 => (x"81",x"c8",x"49",x"6a"),
  1347 => (x"87",x"fa",x"dd",x"ff"),
  1348 => (x"66",x"d0",x"86",x"c8"),
  1349 => (x"a8",x"b7",x"c0",x"48"),
  1350 => (x"c1",x"87",x"c4",x"01"),
  1351 => (x"d0",x"87",x"c8",x"4d"),
  1352 => (x"88",x"c1",x"48",x"66"),
  1353 => (x"d4",x"58",x"a6",x"d4"),
  1354 => (x"f4",x"ca",x"02",x"66"),
  1355 => (x"66",x"c0",x"c1",x"87"),
  1356 => (x"ca",x"03",x"ad",x"b7"),
  1357 => (x"d4",x"ff",x"87",x"eb"),
  1358 => (x"78",x"ff",x"c3",x"48"),
  1359 => (x"ff",x"48",x"a6",x"d4"),
  1360 => (x"d4",x"78",x"bf",x"d4"),
  1361 => (x"c6",x"c1",x"48",x"66"),
  1362 => (x"58",x"a6",x"c4",x"88"),
  1363 => (x"c0",x"02",x"98",x"70"),
  1364 => (x"c9",x"48",x"87",x"e6"),
  1365 => (x"58",x"a6",x"c4",x"88"),
  1366 => (x"c4",x"02",x"98",x"70"),
  1367 => (x"c1",x"48",x"87",x"d5"),
  1368 => (x"58",x"a6",x"c4",x"88"),
  1369 => (x"c1",x"02",x"98",x"70"),
  1370 => (x"c4",x"48",x"87",x"e3"),
  1371 => (x"70",x"58",x"a6",x"88"),
  1372 => (x"fe",x"c3",x"02",x"98"),
  1373 => (x"87",x"d3",x"c9",x"87"),
  1374 => (x"c1",x"05",x"66",x"d8"),
  1375 => (x"d4",x"ff",x"87",x"c5"),
  1376 => (x"78",x"ff",x"c3",x"48"),
  1377 => (x"1e",x"ca",x"1e",x"c0"),
  1378 => (x"93",x"cc",x"4b",x"75"),
  1379 => (x"83",x"66",x"c0",x"c1"),
  1380 => (x"6c",x"4c",x"a3",x"c4"),
  1381 => (x"f1",x"db",x"ff",x"49"),
  1382 => (x"de",x"1e",x"c1",x"87"),
  1383 => (x"ff",x"49",x"6c",x"1e"),
  1384 => (x"d0",x"87",x"e7",x"db"),
  1385 => (x"49",x"a3",x"c8",x"86"),
  1386 => (x"79",x"c0",x"cc",x"c1"),
  1387 => (x"ad",x"b7",x"66",x"d0"),
  1388 => (x"c1",x"87",x"c5",x"04"),
  1389 => (x"87",x"da",x"c8",x"85"),
  1390 => (x"c1",x"48",x"66",x"d0"),
  1391 => (x"58",x"a6",x"d4",x"88"),
  1392 => (x"ff",x"87",x"cf",x"c8"),
  1393 => (x"d8",x"87",x"ec",x"da"),
  1394 => (x"c5",x"c8",x"58",x"a6"),
  1395 => (x"f3",x"dc",x"ff",x"87"),
  1396 => (x"58",x"a6",x"cc",x"87"),
  1397 => (x"a8",x"b7",x"66",x"cc"),
  1398 => (x"cc",x"87",x"c6",x"06"),
  1399 => (x"66",x"c8",x"48",x"a6"),
  1400 => (x"df",x"dc",x"ff",x"78"),
  1401 => (x"a8",x"ec",x"c0",x"87"),
  1402 => (x"87",x"c7",x"c2",x"05"),
  1403 => (x"c1",x"05",x"66",x"d8"),
  1404 => (x"49",x"75",x"87",x"f7"),
  1405 => (x"f8",x"c0",x"91",x"cc"),
  1406 => (x"a1",x"c4",x"81",x"66"),
  1407 => (x"c1",x"4c",x"6a",x"4a"),
  1408 => (x"66",x"c8",x"4a",x"a1"),
  1409 => (x"79",x"97",x"c2",x"52"),
  1410 => (x"cc",x"c1",x"81",x"c8"),
  1411 => (x"d4",x"ff",x"79",x"ce"),
  1412 => (x"78",x"ff",x"c3",x"48"),
  1413 => (x"ff",x"48",x"a6",x"d4"),
  1414 => (x"d4",x"78",x"bf",x"d4"),
  1415 => (x"e8",x"c0",x"02",x"66"),
  1416 => (x"fb",x"c0",x"48",x"87"),
  1417 => (x"e0",x"c0",x"02",x"a8"),
  1418 => (x"97",x"66",x"d4",x"87"),
  1419 => (x"ff",x"84",x"c1",x"7c"),
  1420 => (x"ff",x"c3",x"48",x"d4"),
  1421 => (x"48",x"a6",x"d4",x"78"),
  1422 => (x"78",x"bf",x"d4",x"ff"),
  1423 => (x"c8",x"02",x"66",x"d4"),
  1424 => (x"fb",x"c0",x"48",x"87"),
  1425 => (x"e0",x"ff",x"05",x"a8"),
  1426 => (x"54",x"e0",x"c0",x"87"),
  1427 => (x"c0",x"54",x"c1",x"c2"),
  1428 => (x"66",x"d0",x"7c",x"97"),
  1429 => (x"c5",x"04",x"ad",x"b7"),
  1430 => (x"c5",x"85",x"c1",x"87"),
  1431 => (x"66",x"d0",x"87",x"f4"),
  1432 => (x"d4",x"88",x"c1",x"48"),
  1433 => (x"e9",x"c5",x"58",x"a6"),
  1434 => (x"c6",x"d8",x"ff",x"87"),
  1435 => (x"58",x"a6",x"d8",x"87"),
  1436 => (x"c8",x"87",x"df",x"c5"),
  1437 => (x"66",x"d8",x"48",x"66"),
  1438 => (x"c4",x"c5",x"05",x"a8"),
  1439 => (x"48",x"a6",x"dc",x"87"),
  1440 => (x"d9",x"ff",x"78",x"c0"),
  1441 => (x"a6",x"d8",x"87",x"fe"),
  1442 => (x"f7",x"d9",x"ff",x"58"),
  1443 => (x"a6",x"e4",x"c0",x"87"),
  1444 => (x"a8",x"ec",x"c0",x"58"),
  1445 => (x"87",x"ca",x"c0",x"05"),
  1446 => (x"48",x"a6",x"e0",x"c0"),
  1447 => (x"c0",x"78",x"66",x"d4"),
  1448 => (x"d4",x"ff",x"87",x"c6"),
  1449 => (x"78",x"ff",x"c3",x"48"),
  1450 => (x"91",x"cc",x"49",x"75"),
  1451 => (x"48",x"66",x"f8",x"c0"),
  1452 => (x"a6",x"c4",x"80",x"71"),
  1453 => (x"c3",x"49",x"6e",x"58"),
  1454 => (x"51",x"66",x"d4",x"81"),
  1455 => (x"49",x"66",x"e0",x"c0"),
  1456 => (x"66",x"d4",x"81",x"c1"),
  1457 => (x"71",x"48",x"c1",x"89"),
  1458 => (x"c1",x"49",x"70",x"30"),
  1459 => (x"c1",x"4a",x"6e",x"89"),
  1460 => (x"97",x"09",x"72",x"82"),
  1461 => (x"48",x"6e",x"09",x"79"),
  1462 => (x"e5",x"c2",x"50",x"c2"),
  1463 => (x"d4",x"49",x"bf",x"d0"),
  1464 => (x"97",x"29",x"b7",x"66"),
  1465 => (x"71",x"48",x"4a",x"6a"),
  1466 => (x"a6",x"e8",x"c0",x"98"),
  1467 => (x"c4",x"48",x"6e",x"58"),
  1468 => (x"58",x"a6",x"c8",x"80"),
  1469 => (x"4c",x"bf",x"66",x"c4"),
  1470 => (x"c8",x"48",x"66",x"d8"),
  1471 => (x"c0",x"02",x"a8",x"66"),
  1472 => (x"e0",x"c0",x"87",x"c9"),
  1473 => (x"78",x"c0",x"48",x"a6"),
  1474 => (x"c0",x"87",x"c6",x"c0"),
  1475 => (x"c1",x"48",x"a6",x"e0"),
  1476 => (x"66",x"e0",x"c0",x"78"),
  1477 => (x"1e",x"e0",x"c0",x"1e"),
  1478 => (x"d5",x"ff",x"49",x"74"),
  1479 => (x"86",x"c8",x"87",x"ec"),
  1480 => (x"c0",x"58",x"a6",x"d8"),
  1481 => (x"c1",x"06",x"a8",x"b7"),
  1482 => (x"66",x"d4",x"87",x"da"),
  1483 => (x"bf",x"66",x"c4",x"84"),
  1484 => (x"81",x"e0",x"c0",x"49"),
  1485 => (x"c1",x"4b",x"89",x"74"),
  1486 => (x"71",x"4a",x"f2",x"c2"),
  1487 => (x"87",x"e0",x"e5",x"fe"),
  1488 => (x"66",x"dc",x"84",x"c2"),
  1489 => (x"c0",x"80",x"c1",x"48"),
  1490 => (x"c0",x"58",x"a6",x"e0"),
  1491 => (x"c1",x"49",x"66",x"e4"),
  1492 => (x"02",x"a9",x"70",x"81"),
  1493 => (x"c0",x"87",x"c9",x"c0"),
  1494 => (x"c0",x"48",x"a6",x"e0"),
  1495 => (x"87",x"c6",x"c0",x"78"),
  1496 => (x"48",x"a6",x"e0",x"c0"),
  1497 => (x"e0",x"c0",x"78",x"c1"),
  1498 => (x"66",x"c8",x"1e",x"66"),
  1499 => (x"e0",x"c0",x"49",x"bf"),
  1500 => (x"71",x"89",x"74",x"81"),
  1501 => (x"ff",x"49",x"74",x"1e"),
  1502 => (x"c8",x"87",x"cf",x"d4"),
  1503 => (x"a8",x"b7",x"c0",x"86"),
  1504 => (x"87",x"fe",x"fe",x"01"),
  1505 => (x"c0",x"02",x"66",x"dc"),
  1506 => (x"49",x"6e",x"87",x"d2"),
  1507 => (x"66",x"dc",x"81",x"c2"),
  1508 => (x"c8",x"49",x"6e",x"51"),
  1509 => (x"ef",x"cc",x"c1",x"81"),
  1510 => (x"87",x"cd",x"c0",x"79"),
  1511 => (x"81",x"c2",x"49",x"6e"),
  1512 => (x"c8",x"49",x"6e",x"51"),
  1513 => (x"d5",x"d0",x"c1",x"81"),
  1514 => (x"b7",x"66",x"d0",x"79"),
  1515 => (x"c5",x"c0",x"04",x"ad"),
  1516 => (x"c0",x"85",x"c1",x"87"),
  1517 => (x"66",x"d0",x"87",x"dc"),
  1518 => (x"d4",x"88",x"c1",x"48"),
  1519 => (x"d1",x"c0",x"58",x"a6"),
  1520 => (x"ee",x"d2",x"ff",x"87"),
  1521 => (x"58",x"a6",x"d8",x"87"),
  1522 => (x"ff",x"87",x"c7",x"c0"),
  1523 => (x"d8",x"87",x"e4",x"d2"),
  1524 => (x"66",x"d4",x"58",x"a6"),
  1525 => (x"87",x"c9",x"c0",x"02"),
  1526 => (x"b7",x"66",x"c0",x"c1"),
  1527 => (x"d5",x"f5",x"04",x"ad"),
  1528 => (x"ad",x"b7",x"c7",x"87"),
  1529 => (x"87",x"dc",x"c0",x"03"),
  1530 => (x"91",x"cc",x"49",x"75"),
  1531 => (x"81",x"66",x"f8",x"c0"),
  1532 => (x"6a",x"4a",x"a1",x"c4"),
  1533 => (x"c8",x"52",x"c0",x"4a"),
  1534 => (x"c1",x"79",x"c0",x"81"),
  1535 => (x"ad",x"b7",x"c7",x"85"),
  1536 => (x"87",x"e4",x"ff",x"04"),
  1537 => (x"c0",x"02",x"66",x"d8"),
  1538 => (x"f8",x"c0",x"87",x"eb"),
  1539 => (x"d4",x"c1",x"49",x"66"),
  1540 => (x"66",x"f8",x"c0",x"81"),
  1541 => (x"82",x"d5",x"c1",x"4a"),
  1542 => (x"51",x"c2",x"52",x"c0"),
  1543 => (x"49",x"66",x"f8",x"c0"),
  1544 => (x"c1",x"81",x"dc",x"c1"),
  1545 => (x"c0",x"79",x"ce",x"cc"),
  1546 => (x"c1",x"49",x"66",x"f8"),
  1547 => (x"c2",x"c1",x"81",x"d8"),
  1548 => (x"d6",x"c0",x"79",x"f5"),
  1549 => (x"66",x"f8",x"c0",x"87"),
  1550 => (x"81",x"d8",x"c1",x"49"),
  1551 => (x"79",x"fc",x"c2",x"c1"),
  1552 => (x"49",x"66",x"f8",x"c0"),
  1553 => (x"c2",x"81",x"dc",x"c1"),
  1554 => (x"c1",x"79",x"e5",x"ca"),
  1555 => (x"c0",x"4a",x"e6",x"d0"),
  1556 => (x"c1",x"49",x"66",x"f8"),
  1557 => (x"79",x"72",x"81",x"e8"),
  1558 => (x"48",x"bf",x"d0",x"ff"),
  1559 => (x"98",x"c0",x"c0",x"c8"),
  1560 => (x"70",x"58",x"a6",x"c4"),
  1561 => (x"d1",x"c0",x"02",x"98"),
  1562 => (x"bf",x"d0",x"ff",x"87"),
  1563 => (x"c0",x"c0",x"c8",x"48"),
  1564 => (x"58",x"a6",x"c4",x"98"),
  1565 => (x"ff",x"05",x"98",x"70"),
  1566 => (x"d0",x"ff",x"87",x"ef"),
  1567 => (x"78",x"e0",x"c0",x"48"),
  1568 => (x"ff",x"48",x"66",x"cc"),
  1569 => (x"d1",x"ff",x"8e",x"d8"),
  1570 => (x"c7",x"1e",x"87",x"f2"),
  1571 => (x"c1",x"1e",x"c0",x"1e"),
  1572 => (x"c2",x"1e",x"d0",x"e4"),
  1573 => (x"49",x"bf",x"d4",x"e5"),
  1574 => (x"c1",x"87",x"d0",x"ef"),
  1575 => (x"c0",x"49",x"d0",x"e4"),
  1576 => (x"f4",x"87",x"e2",x"e7"),
  1577 => (x"1e",x"4f",x"26",x"8e"),
  1578 => (x"c2",x"87",x"c6",x"ca"),
  1579 => (x"c0",x"48",x"f0",x"e5"),
  1580 => (x"48",x"d4",x"ff",x"50"),
  1581 => (x"c1",x"78",x"ff",x"c3"),
  1582 => (x"fe",x"49",x"c3",x"c3"),
  1583 => (x"fe",x"87",x"fd",x"de"),
  1584 => (x"70",x"87",x"c8",x"e8"),
  1585 => (x"87",x"cd",x"02",x"98"),
  1586 => (x"87",x"c5",x"f4",x"fe"),
  1587 => (x"c4",x"02",x"98",x"70"),
  1588 => (x"c2",x"4a",x"c1",x"87"),
  1589 => (x"72",x"4a",x"c0",x"87"),
  1590 => (x"87",x"c8",x"02",x"9a"),
  1591 => (x"49",x"cd",x"c3",x"c1"),
  1592 => (x"87",x"d8",x"de",x"fe"),
  1593 => (x"bf",x"c0",x"d7",x"c2"),
  1594 => (x"e3",x"d5",x"ff",x"49"),
  1595 => (x"e8",x"e5",x"c2",x"87"),
  1596 => (x"c2",x"78",x"c0",x"48"),
  1597 => (x"c0",x"48",x"d4",x"e5"),
  1598 => (x"cd",x"fe",x"49",x"78"),
  1599 => (x"87",x"dd",x"c3",x"87"),
  1600 => (x"c0",x"87",x"c2",x"c9"),
  1601 => (x"ff",x"87",x"ed",x"e6"),
  1602 => (x"4f",x"26",x"87",x"f6"),
  1603 => (x"00",x"00",x"10",x"d0"),
  1604 => (x"00",x"00",x"00",x"02"),
  1605 => (x"00",x"00",x"29",x"80"),
  1606 => (x"00",x"00",x"10",x"32"),
  1607 => (x"00",x"00",x"00",x"02"),
  1608 => (x"00",x"00",x"29",x"9e"),
  1609 => (x"00",x"00",x"10",x"32"),
  1610 => (x"00",x"00",x"00",x"02"),
  1611 => (x"00",x"00",x"29",x"bc"),
  1612 => (x"00",x"00",x"10",x"32"),
  1613 => (x"00",x"00",x"00",x"02"),
  1614 => (x"00",x"00",x"29",x"da"),
  1615 => (x"00",x"00",x"10",x"32"),
  1616 => (x"00",x"00",x"00",x"02"),
  1617 => (x"00",x"00",x"29",x"f8"),
  1618 => (x"00",x"00",x"10",x"32"),
  1619 => (x"00",x"00",x"00",x"02"),
  1620 => (x"00",x"00",x"2a",x"16"),
  1621 => (x"00",x"00",x"10",x"32"),
  1622 => (x"00",x"00",x"00",x"02"),
  1623 => (x"00",x"00",x"2a",x"34"),
  1624 => (x"00",x"00",x"10",x"32"),
  1625 => (x"00",x"00",x"00",x"02"),
  1626 => (x"00",x"00",x"00",x"00"),
  1627 => (x"00",x"00",x"13",x"0e"),
  1628 => (x"00",x"00",x"00",x"00"),
  1629 => (x"00",x"00",x"00",x"00"),
  1630 => (x"00",x"00",x"11",x"02"),
  1631 => (x"d5",x"c1",x"1e",x"1e"),
  1632 => (x"58",x"a6",x"c4",x"87"),
  1633 => (x"1e",x"4f",x"26",x"26"),
  1634 => (x"f0",x"fe",x"4a",x"71"),
  1635 => (x"cd",x"78",x"c0",x"48"),
  1636 => (x"c1",x"0a",x"7a",x"0a"),
  1637 => (x"fe",x"49",x"dd",x"e6"),
  1638 => (x"26",x"87",x"e1",x"db"),
  1639 => (x"74",x"65",x"53",x"4f"),
  1640 => (x"6e",x"61",x"68",x"20"),
  1641 => (x"72",x"65",x"6c",x"64"),
  1642 => (x"6e",x"49",x"00",x"0a"),
  1643 => (x"74",x"6e",x"69",x"20"),
  1644 => (x"75",x"72",x"72",x"65"),
  1645 => (x"63",x"20",x"74",x"70"),
  1646 => (x"74",x"73",x"6e",x"6f"),
  1647 => (x"74",x"63",x"75",x"72"),
  1648 => (x"00",x"0a",x"72",x"6f"),
  1649 => (x"ea",x"e6",x"c1",x"1e"),
  1650 => (x"ef",x"da",x"fe",x"49"),
  1651 => (x"fc",x"e5",x"c1",x"87"),
  1652 => (x"87",x"f3",x"fe",x"49"),
  1653 => (x"fe",x"1e",x"4f",x"26"),
  1654 => (x"26",x"48",x"bf",x"f0"),
  1655 => (x"f0",x"fe",x"1e",x"4f"),
  1656 => (x"26",x"78",x"c1",x"48"),
  1657 => (x"f0",x"fe",x"1e",x"4f"),
  1658 => (x"26",x"78",x"c0",x"48"),
  1659 => (x"4a",x"71",x"1e",x"4f"),
  1660 => (x"a2",x"c4",x"7a",x"c0"),
  1661 => (x"c8",x"79",x"c0",x"49"),
  1662 => (x"79",x"c0",x"49",x"a2"),
  1663 => (x"c0",x"49",x"a2",x"cc"),
  1664 => (x"0e",x"4f",x"26",x"79"),
  1665 => (x"0e",x"5c",x"5b",x"5e"),
  1666 => (x"4c",x"71",x"86",x"f8"),
  1667 => (x"cc",x"49",x"a4",x"c8"),
  1668 => (x"48",x"6b",x"4b",x"a4"),
  1669 => (x"a6",x"c4",x"80",x"c1"),
  1670 => (x"c8",x"98",x"cf",x"58"),
  1671 => (x"48",x"69",x"58",x"a6"),
  1672 => (x"05",x"a8",x"66",x"c4"),
  1673 => (x"48",x"6b",x"87",x"d4"),
  1674 => (x"a6",x"c4",x"80",x"c1"),
  1675 => (x"c8",x"98",x"cf",x"58"),
  1676 => (x"48",x"69",x"58",x"a6"),
  1677 => (x"02",x"a8",x"66",x"c4"),
  1678 => (x"e8",x"fe",x"87",x"ec"),
  1679 => (x"a4",x"d0",x"c1",x"87"),
  1680 => (x"c4",x"48",x"6b",x"49"),
  1681 => (x"58",x"a6",x"c4",x"90"),
  1682 => (x"66",x"d4",x"81",x"70"),
  1683 => (x"c1",x"48",x"6b",x"79"),
  1684 => (x"58",x"a6",x"c8",x"80"),
  1685 => (x"7b",x"70",x"98",x"cf"),
  1686 => (x"fd",x"87",x"d2",x"c1"),
  1687 => (x"8e",x"f8",x"87",x"ff"),
  1688 => (x"4d",x"26",x"87",x"c2"),
  1689 => (x"4b",x"26",x"4c",x"26"),
  1690 => (x"5e",x"0e",x"4f",x"26"),
  1691 => (x"0e",x"5d",x"5c",x"5b"),
  1692 => (x"4d",x"71",x"86",x"f8"),
  1693 => (x"6d",x"4c",x"a5",x"c4"),
  1694 => (x"05",x"a8",x"6c",x"48"),
  1695 => (x"48",x"ff",x"87",x"c5"),
  1696 => (x"fd",x"87",x"e5",x"c0"),
  1697 => (x"a5",x"d0",x"87",x"df"),
  1698 => (x"c4",x"48",x"6c",x"4b"),
  1699 => (x"58",x"a6",x"c4",x"90"),
  1700 => (x"4b",x"6b",x"83",x"70"),
  1701 => (x"6c",x"9b",x"ff",x"c3"),
  1702 => (x"c8",x"80",x"c1",x"48"),
  1703 => (x"98",x"cf",x"58",x"a6"),
  1704 => (x"f8",x"fc",x"7c",x"70"),
  1705 => (x"48",x"49",x"73",x"87"),
  1706 => (x"f5",x"fe",x"8e",x"f8"),
  1707 => (x"1e",x"73",x"1e",x"87"),
  1708 => (x"f0",x"fc",x"86",x"f8"),
  1709 => (x"4b",x"bf",x"e0",x"87"),
  1710 => (x"c0",x"e0",x"c0",x"49"),
  1711 => (x"e7",x"c0",x"02",x"99"),
  1712 => (x"c3",x"4a",x"73",x"87"),
  1713 => (x"e9",x"c2",x"9a",x"ff"),
  1714 => (x"c4",x"48",x"bf",x"d2"),
  1715 => (x"58",x"a6",x"c4",x"90"),
  1716 => (x"49",x"e2",x"e9",x"c2"),
  1717 => (x"79",x"72",x"81",x"70"),
  1718 => (x"bf",x"d2",x"e9",x"c2"),
  1719 => (x"c8",x"80",x"c1",x"48"),
  1720 => (x"98",x"cf",x"58",x"a6"),
  1721 => (x"58",x"d6",x"e9",x"c2"),
  1722 => (x"c0",x"d0",x"49",x"73"),
  1723 => (x"f2",x"c0",x"02",x"99"),
  1724 => (x"da",x"e9",x"c2",x"87"),
  1725 => (x"e9",x"c2",x"48",x"bf"),
  1726 => (x"02",x"a8",x"bf",x"de"),
  1727 => (x"c2",x"87",x"e4",x"c0"),
  1728 => (x"48",x"bf",x"da",x"e9"),
  1729 => (x"a6",x"c4",x"90",x"c4"),
  1730 => (x"e2",x"ea",x"c2",x"58"),
  1731 => (x"e0",x"81",x"70",x"49"),
  1732 => (x"c2",x"78",x"69",x"48"),
  1733 => (x"48",x"bf",x"da",x"e9"),
  1734 => (x"a6",x"c8",x"80",x"c1"),
  1735 => (x"c2",x"98",x"cf",x"58"),
  1736 => (x"fa",x"58",x"de",x"e9"),
  1737 => (x"a6",x"c4",x"87",x"f0"),
  1738 => (x"87",x"f1",x"fa",x"58"),
  1739 => (x"f5",x"fc",x"8e",x"f8"),
  1740 => (x"e9",x"c2",x"1e",x"87"),
  1741 => (x"f4",x"fa",x"49",x"d2"),
  1742 => (x"ed",x"ea",x"c1",x"87"),
  1743 => (x"87",x"c7",x"f9",x"49"),
  1744 => (x"26",x"87",x"f5",x"c3"),
  1745 => (x"1e",x"73",x"1e",x"4f"),
  1746 => (x"49",x"d2",x"e9",x"c2"),
  1747 => (x"70",x"87",x"db",x"fc"),
  1748 => (x"aa",x"b7",x"c0",x"4a"),
  1749 => (x"87",x"cc",x"c2",x"04"),
  1750 => (x"05",x"aa",x"f0",x"c3"),
  1751 => (x"ef",x"c1",x"87",x"c9"),
  1752 => (x"78",x"c1",x"48",x"f0"),
  1753 => (x"c3",x"87",x"ed",x"c1"),
  1754 => (x"c9",x"05",x"aa",x"e0"),
  1755 => (x"f4",x"ef",x"c1",x"87"),
  1756 => (x"c1",x"78",x"c1",x"48"),
  1757 => (x"ef",x"c1",x"87",x"de"),
  1758 => (x"c6",x"02",x"bf",x"f4"),
  1759 => (x"a2",x"c0",x"c2",x"87"),
  1760 => (x"72",x"87",x"c2",x"4b"),
  1761 => (x"f0",x"ef",x"c1",x"4b"),
  1762 => (x"e0",x"c0",x"02",x"bf"),
  1763 => (x"c4",x"49",x"73",x"87"),
  1764 => (x"c1",x"91",x"29",x"b7"),
  1765 => (x"73",x"81",x"f8",x"ef"),
  1766 => (x"c2",x"9a",x"cf",x"4a"),
  1767 => (x"72",x"48",x"c1",x"92"),
  1768 => (x"ff",x"4a",x"70",x"30"),
  1769 => (x"69",x"48",x"72",x"ba"),
  1770 => (x"db",x"79",x"70",x"98"),
  1771 => (x"c4",x"49",x"73",x"87"),
  1772 => (x"c1",x"91",x"29",x"b7"),
  1773 => (x"73",x"81",x"f8",x"ef"),
  1774 => (x"c2",x"9a",x"cf",x"4a"),
  1775 => (x"72",x"48",x"c3",x"92"),
  1776 => (x"48",x"4a",x"70",x"30"),
  1777 => (x"79",x"70",x"b0",x"69"),
  1778 => (x"48",x"f4",x"ef",x"c1"),
  1779 => (x"ef",x"c1",x"78",x"c0"),
  1780 => (x"78",x"c0",x"48",x"f0"),
  1781 => (x"49",x"d2",x"e9",x"c2"),
  1782 => (x"70",x"87",x"cf",x"fa"),
  1783 => (x"aa",x"b7",x"c0",x"4a"),
  1784 => (x"87",x"f4",x"fd",x"03"),
  1785 => (x"87",x"c4",x"48",x"c0"),
  1786 => (x"4c",x"26",x"4d",x"26"),
  1787 => (x"4f",x"26",x"4b",x"26"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"72",x"4a",x"c0",x"1e"),
  1807 => (x"c1",x"91",x"c4",x"49"),
  1808 => (x"c0",x"81",x"f8",x"ef"),
  1809 => (x"d0",x"82",x"c1",x"79"),
  1810 => (x"ee",x"04",x"aa",x"b7"),
  1811 => (x"0e",x"4f",x"26",x"87"),
  1812 => (x"5d",x"5c",x"5b",x"5e"),
  1813 => (x"f6",x"4d",x"71",x"0e"),
  1814 => (x"4a",x"75",x"87",x"cb"),
  1815 => (x"92",x"2a",x"b7",x"c4"),
  1816 => (x"82",x"f8",x"ef",x"c1"),
  1817 => (x"9c",x"cf",x"4c",x"75"),
  1818 => (x"49",x"6a",x"94",x"c2"),
  1819 => (x"c3",x"2b",x"74",x"4b"),
  1820 => (x"74",x"48",x"c2",x"9b"),
  1821 => (x"ff",x"4c",x"70",x"30"),
  1822 => (x"71",x"48",x"74",x"bc"),
  1823 => (x"f5",x"7a",x"70",x"98"),
  1824 => (x"48",x"73",x"87",x"db"),
  1825 => (x"1e",x"87",x"e1",x"fd"),
  1826 => (x"bf",x"d0",x"ff",x"1e"),
  1827 => (x"c0",x"c0",x"c8",x"48"),
  1828 => (x"58",x"a6",x"c4",x"98"),
  1829 => (x"d0",x"02",x"98",x"70"),
  1830 => (x"bf",x"d0",x"ff",x"87"),
  1831 => (x"c0",x"c0",x"c8",x"48"),
  1832 => (x"58",x"a6",x"c4",x"98"),
  1833 => (x"f0",x"05",x"98",x"70"),
  1834 => (x"48",x"d0",x"ff",x"87"),
  1835 => (x"71",x"78",x"e1",x"c4"),
  1836 => (x"08",x"d4",x"ff",x"48"),
  1837 => (x"48",x"66",x"c8",x"78"),
  1838 => (x"78",x"08",x"d4",x"ff"),
  1839 => (x"1e",x"4f",x"26",x"26"),
  1840 => (x"c8",x"4a",x"71",x"1e"),
  1841 => (x"72",x"1e",x"49",x"66"),
  1842 => (x"87",x"fb",x"fe",x"49"),
  1843 => (x"d0",x"ff",x"86",x"c4"),
  1844 => (x"c0",x"c8",x"48",x"bf"),
  1845 => (x"a6",x"c4",x"98",x"c0"),
  1846 => (x"02",x"98",x"70",x"58"),
  1847 => (x"d0",x"ff",x"87",x"d0"),
  1848 => (x"c0",x"c8",x"48",x"bf"),
  1849 => (x"a6",x"c4",x"98",x"c0"),
  1850 => (x"05",x"98",x"70",x"58"),
  1851 => (x"d0",x"ff",x"87",x"f0"),
  1852 => (x"78",x"e0",x"c0",x"48"),
  1853 => (x"1e",x"4f",x"26",x"26"),
  1854 => (x"4b",x"71",x"1e",x"73"),
  1855 => (x"73",x"1e",x"66",x"c8"),
  1856 => (x"a2",x"e0",x"c1",x"4a"),
  1857 => (x"87",x"f7",x"fe",x"49"),
  1858 => (x"26",x"87",x"c4",x"26"),
  1859 => (x"26",x"4c",x"26",x"4d"),
  1860 => (x"1e",x"4f",x"26",x"4b"),
  1861 => (x"bf",x"d0",x"ff",x"1e"),
  1862 => (x"c0",x"c0",x"c8",x"48"),
  1863 => (x"58",x"a6",x"c4",x"98"),
  1864 => (x"d0",x"02",x"98",x"70"),
  1865 => (x"bf",x"d0",x"ff",x"87"),
  1866 => (x"c0",x"c0",x"c8",x"48"),
  1867 => (x"58",x"a6",x"c4",x"98"),
  1868 => (x"f0",x"05",x"98",x"70"),
  1869 => (x"48",x"d0",x"ff",x"87"),
  1870 => (x"71",x"78",x"c9",x"c4"),
  1871 => (x"08",x"d4",x"ff",x"48"),
  1872 => (x"4f",x"26",x"26",x"78"),
  1873 => (x"4a",x"71",x"1e",x"1e"),
  1874 => (x"87",x"c7",x"ff",x"49"),
  1875 => (x"48",x"bf",x"d0",x"ff"),
  1876 => (x"98",x"c0",x"c0",x"c8"),
  1877 => (x"70",x"58",x"a6",x"c4"),
  1878 => (x"87",x"d0",x"02",x"98"),
  1879 => (x"48",x"bf",x"d0",x"ff"),
  1880 => (x"98",x"c0",x"c0",x"c8"),
  1881 => (x"70",x"58",x"a6",x"c4"),
  1882 => (x"87",x"f0",x"05",x"98"),
  1883 => (x"c8",x"48",x"d0",x"ff"),
  1884 => (x"4f",x"26",x"26",x"78"),
  1885 => (x"1e",x"1e",x"73",x"1e"),
  1886 => (x"eb",x"c2",x"4b",x"71"),
  1887 => (x"c3",x"02",x"bf",x"ee"),
  1888 => (x"87",x"cc",x"c3",x"87"),
  1889 => (x"48",x"bf",x"d0",x"ff"),
  1890 => (x"98",x"c0",x"c0",x"c8"),
  1891 => (x"70",x"58",x"a6",x"c4"),
  1892 => (x"87",x"d0",x"02",x"98"),
  1893 => (x"48",x"bf",x"d0",x"ff"),
  1894 => (x"98",x"c0",x"c0",x"c8"),
  1895 => (x"70",x"58",x"a6",x"c4"),
  1896 => (x"87",x"f0",x"05",x"98"),
  1897 => (x"c4",x"48",x"d0",x"ff"),
  1898 => (x"48",x"73",x"78",x"c9"),
  1899 => (x"ff",x"b0",x"e0",x"c0"),
  1900 => (x"c2",x"78",x"08",x"d4"),
  1901 => (x"c0",x"48",x"e2",x"eb"),
  1902 => (x"02",x"66",x"cc",x"78"),
  1903 => (x"ff",x"c3",x"87",x"c5"),
  1904 => (x"c0",x"87",x"c2",x"49"),
  1905 => (x"ea",x"eb",x"c2",x"49"),
  1906 => (x"02",x"66",x"d0",x"59"),
  1907 => (x"d5",x"c5",x"87",x"c6"),
  1908 => (x"87",x"c4",x"4a",x"d5"),
  1909 => (x"4a",x"ff",x"ff",x"cf"),
  1910 => (x"5a",x"ee",x"eb",x"c2"),
  1911 => (x"48",x"ee",x"eb",x"c2"),
  1912 => (x"c4",x"26",x"78",x"c1"),
  1913 => (x"26",x"4d",x"26",x"87"),
  1914 => (x"26",x"4b",x"26",x"4c"),
  1915 => (x"5b",x"5e",x"0e",x"4f"),
  1916 => (x"71",x"0e",x"5d",x"5c"),
  1917 => (x"ea",x"eb",x"c2",x"4a"),
  1918 => (x"9a",x"72",x"4c",x"bf"),
  1919 => (x"49",x"87",x"cb",x"02"),
  1920 => (x"f6",x"c1",x"91",x"c8"),
  1921 => (x"83",x"71",x"4b",x"ee"),
  1922 => (x"fa",x"c1",x"87",x"c4"),
  1923 => (x"4d",x"c0",x"4b",x"ee"),
  1924 => (x"99",x"74",x"49",x"13"),
  1925 => (x"bf",x"e6",x"eb",x"c2"),
  1926 => (x"ff",x"b8",x"71",x"48"),
  1927 => (x"c1",x"78",x"08",x"d4"),
  1928 => (x"c8",x"85",x"2c",x"b7"),
  1929 => (x"e7",x"04",x"ad",x"b7"),
  1930 => (x"e2",x"eb",x"c2",x"87"),
  1931 => (x"80",x"c8",x"48",x"bf"),
  1932 => (x"58",x"e6",x"eb",x"c2"),
  1933 => (x"1e",x"87",x"ee",x"fe"),
  1934 => (x"4b",x"71",x"1e",x"73"),
  1935 => (x"02",x"9a",x"4a",x"13"),
  1936 => (x"49",x"72",x"87",x"cb"),
  1937 => (x"13",x"87",x"e6",x"fe"),
  1938 => (x"f5",x"05",x"9a",x"4a"),
  1939 => (x"87",x"d9",x"fe",x"87"),
  1940 => (x"eb",x"c2",x"1e",x"1e"),
  1941 => (x"c2",x"49",x"bf",x"e2"),
  1942 => (x"c1",x"48",x"e2",x"eb"),
  1943 => (x"c0",x"c4",x"78",x"a1"),
  1944 => (x"db",x"03",x"a9",x"b7"),
  1945 => (x"48",x"d4",x"ff",x"87"),
  1946 => (x"bf",x"e6",x"eb",x"c2"),
  1947 => (x"e2",x"eb",x"c2",x"78"),
  1948 => (x"eb",x"c2",x"49",x"bf"),
  1949 => (x"a1",x"c1",x"48",x"e2"),
  1950 => (x"b7",x"c0",x"c4",x"78"),
  1951 => (x"87",x"e5",x"04",x"a9"),
  1952 => (x"48",x"bf",x"d0",x"ff"),
  1953 => (x"98",x"c0",x"c0",x"c8"),
  1954 => (x"70",x"58",x"a6",x"c4"),
  1955 => (x"87",x"d0",x"02",x"98"),
  1956 => (x"48",x"bf",x"d0",x"ff"),
  1957 => (x"98",x"c0",x"c0",x"c8"),
  1958 => (x"70",x"58",x"a6",x"c4"),
  1959 => (x"87",x"f0",x"05",x"98"),
  1960 => (x"c8",x"48",x"d0",x"ff"),
  1961 => (x"ee",x"eb",x"c2",x"78"),
  1962 => (x"26",x"78",x"c0",x"48"),
  1963 => (x"00",x"00",x"4f",x"26"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"5f",x"5f",x"00"),
  1967 => (x"03",x"00",x"00",x"00"),
  1968 => (x"03",x"03",x"00",x"03"),
  1969 => (x"7f",x"14",x"00",x"00"),
  1970 => (x"7f",x"7f",x"14",x"7f"),
  1971 => (x"24",x"00",x"00",x"14"),
  1972 => (x"3a",x"6b",x"6b",x"2e"),
  1973 => (x"6a",x"4c",x"00",x"12"),
  1974 => (x"56",x"6c",x"18",x"36"),
  1975 => (x"7e",x"30",x"00",x"32"),
  1976 => (x"3a",x"77",x"59",x"4f"),
  1977 => (x"00",x"00",x"40",x"68"),
  1978 => (x"00",x"03",x"07",x"04"),
  1979 => (x"00",x"00",x"00",x"00"),
  1980 => (x"41",x"63",x"3e",x"1c"),
  1981 => (x"00",x"00",x"00",x"00"),
  1982 => (x"1c",x"3e",x"63",x"41"),
  1983 => (x"2a",x"08",x"00",x"00"),
  1984 => (x"3e",x"1c",x"1c",x"3e"),
  1985 => (x"08",x"00",x"08",x"2a"),
  1986 => (x"08",x"3e",x"3e",x"08"),
  1987 => (x"00",x"00",x"00",x"08"),
  1988 => (x"00",x"60",x"e0",x"80"),
  1989 => (x"08",x"00",x"00",x"00"),
  1990 => (x"08",x"08",x"08",x"08"),
  1991 => (x"00",x"00",x"00",x"08"),
  1992 => (x"00",x"60",x"60",x"00"),
  1993 => (x"60",x"40",x"00",x"00"),
  1994 => (x"06",x"0c",x"18",x"30"),
  1995 => (x"3e",x"00",x"01",x"03"),
  1996 => (x"7f",x"4d",x"59",x"7f"),
  1997 => (x"04",x"00",x"00",x"3e"),
  1998 => (x"00",x"7f",x"7f",x"06"),
  1999 => (x"42",x"00",x"00",x"00"),
  2000 => (x"4f",x"59",x"71",x"63"),
  2001 => (x"22",x"00",x"00",x"46"),
  2002 => (x"7f",x"49",x"49",x"63"),
  2003 => (x"1c",x"18",x"00",x"36"),
  2004 => (x"7f",x"7f",x"13",x"16"),
  2005 => (x"27",x"00",x"00",x"10"),
  2006 => (x"7d",x"45",x"45",x"67"),
  2007 => (x"3c",x"00",x"00",x"39"),
  2008 => (x"79",x"49",x"4b",x"7e"),
  2009 => (x"01",x"00",x"00",x"30"),
  2010 => (x"0f",x"79",x"71",x"01"),
  2011 => (x"36",x"00",x"00",x"07"),
  2012 => (x"7f",x"49",x"49",x"7f"),
  2013 => (x"06",x"00",x"00",x"36"),
  2014 => (x"3f",x"69",x"49",x"4f"),
  2015 => (x"00",x"00",x"00",x"1e"),
  2016 => (x"00",x"66",x"66",x"00"),
  2017 => (x"00",x"00",x"00",x"00"),
  2018 => (x"00",x"66",x"e6",x"80"),
  2019 => (x"08",x"00",x"00",x"00"),
  2020 => (x"22",x"14",x"14",x"08"),
  2021 => (x"14",x"00",x"00",x"22"),
  2022 => (x"14",x"14",x"14",x"14"),
  2023 => (x"22",x"00",x"00",x"14"),
  2024 => (x"08",x"14",x"14",x"22"),
  2025 => (x"02",x"00",x"00",x"08"),
  2026 => (x"0f",x"59",x"51",x"03"),
  2027 => (x"7f",x"3e",x"00",x"06"),
  2028 => (x"1f",x"55",x"5d",x"41"),
  2029 => (x"7e",x"00",x"00",x"1e"),
  2030 => (x"7f",x"09",x"09",x"7f"),
  2031 => (x"7f",x"00",x"00",x"7e"),
  2032 => (x"7f",x"49",x"49",x"7f"),
  2033 => (x"1c",x"00",x"00",x"36"),
  2034 => (x"41",x"41",x"63",x"3e"),
  2035 => (x"7f",x"00",x"00",x"41"),
  2036 => (x"3e",x"63",x"41",x"7f"),
  2037 => (x"7f",x"00",x"00",x"1c"),
  2038 => (x"41",x"49",x"49",x"7f"),
  2039 => (x"7f",x"00",x"00",x"41"),
  2040 => (x"01",x"09",x"09",x"7f"),
  2041 => (x"3e",x"00",x"00",x"01"),
  2042 => (x"7b",x"49",x"41",x"7f"),
  2043 => (x"7f",x"00",x"00",x"7a"),
  2044 => (x"7f",x"08",x"08",x"7f"),
  2045 => (x"00",x"00",x"00",x"7f"),
  2046 => (x"41",x"7f",x"7f",x"41"),
  2047 => (x"20",x"00",x"00",x"00"),
  2048 => (x"7f",x"40",x"40",x"60"),
  2049 => (x"7f",x"7f",x"00",x"3f"),
  2050 => (x"63",x"36",x"1c",x"08"),
  2051 => (x"7f",x"00",x"00",x"41"),
  2052 => (x"40",x"40",x"40",x"7f"),
  2053 => (x"7f",x"7f",x"00",x"40"),
  2054 => (x"7f",x"06",x"0c",x"06"),
  2055 => (x"7f",x"7f",x"00",x"7f"),
  2056 => (x"7f",x"18",x"0c",x"06"),
  2057 => (x"3e",x"00",x"00",x"7f"),
  2058 => (x"7f",x"41",x"41",x"7f"),
  2059 => (x"7f",x"00",x"00",x"3e"),
  2060 => (x"0f",x"09",x"09",x"7f"),
  2061 => (x"7f",x"3e",x"00",x"06"),
  2062 => (x"7e",x"7f",x"61",x"41"),
  2063 => (x"7f",x"00",x"00",x"40"),
  2064 => (x"7f",x"19",x"09",x"7f"),
  2065 => (x"26",x"00",x"00",x"66"),
  2066 => (x"7b",x"59",x"4d",x"6f"),
  2067 => (x"01",x"00",x"00",x"32"),
  2068 => (x"01",x"7f",x"7f",x"01"),
  2069 => (x"3f",x"00",x"00",x"01"),
  2070 => (x"7f",x"40",x"40",x"7f"),
  2071 => (x"0f",x"00",x"00",x"3f"),
  2072 => (x"3f",x"70",x"70",x"3f"),
  2073 => (x"7f",x"7f",x"00",x"0f"),
  2074 => (x"7f",x"30",x"18",x"30"),
  2075 => (x"63",x"41",x"00",x"7f"),
  2076 => (x"36",x"1c",x"1c",x"36"),
  2077 => (x"03",x"01",x"41",x"63"),
  2078 => (x"06",x"7c",x"7c",x"06"),
  2079 => (x"71",x"61",x"01",x"03"),
  2080 => (x"43",x"47",x"4d",x"59"),
  2081 => (x"00",x"00",x"00",x"41"),
  2082 => (x"41",x"41",x"7f",x"7f"),
  2083 => (x"03",x"01",x"00",x"00"),
  2084 => (x"30",x"18",x"0c",x"06"),
  2085 => (x"00",x"00",x"40",x"60"),
  2086 => (x"7f",x"7f",x"41",x"41"),
  2087 => (x"0c",x"08",x"00",x"00"),
  2088 => (x"0c",x"06",x"03",x"06"),
  2089 => (x"80",x"80",x"00",x"08"),
  2090 => (x"80",x"80",x"80",x"80"),
  2091 => (x"00",x"00",x"00",x"80"),
  2092 => (x"04",x"07",x"03",x"00"),
  2093 => (x"20",x"00",x"00",x"00"),
  2094 => (x"7c",x"54",x"54",x"74"),
  2095 => (x"7f",x"00",x"00",x"78"),
  2096 => (x"7c",x"44",x"44",x"7f"),
  2097 => (x"38",x"00",x"00",x"38"),
  2098 => (x"44",x"44",x"44",x"7c"),
  2099 => (x"38",x"00",x"00",x"00"),
  2100 => (x"7f",x"44",x"44",x"7c"),
  2101 => (x"38",x"00",x"00",x"7f"),
  2102 => (x"5c",x"54",x"54",x"7c"),
  2103 => (x"04",x"00",x"00",x"18"),
  2104 => (x"05",x"05",x"7f",x"7e"),
  2105 => (x"18",x"00",x"00",x"00"),
  2106 => (x"fc",x"a4",x"a4",x"bc"),
  2107 => (x"7f",x"00",x"00",x"7c"),
  2108 => (x"7c",x"04",x"04",x"7f"),
  2109 => (x"00",x"00",x"00",x"78"),
  2110 => (x"40",x"7d",x"3d",x"00"),
  2111 => (x"80",x"00",x"00",x"00"),
  2112 => (x"7d",x"fd",x"80",x"80"),
  2113 => (x"7f",x"00",x"00",x"00"),
  2114 => (x"6c",x"38",x"10",x"7f"),
  2115 => (x"00",x"00",x"00",x"44"),
  2116 => (x"40",x"7f",x"3f",x"00"),
  2117 => (x"7c",x"7c",x"00",x"00"),
  2118 => (x"7c",x"0c",x"18",x"0c"),
  2119 => (x"7c",x"00",x"00",x"78"),
  2120 => (x"7c",x"04",x"04",x"7c"),
  2121 => (x"38",x"00",x"00",x"78"),
  2122 => (x"7c",x"44",x"44",x"7c"),
  2123 => (x"fc",x"00",x"00",x"38"),
  2124 => (x"3c",x"24",x"24",x"fc"),
  2125 => (x"18",x"00",x"00",x"18"),
  2126 => (x"fc",x"24",x"24",x"3c"),
  2127 => (x"7c",x"00",x"00",x"fc"),
  2128 => (x"0c",x"04",x"04",x"7c"),
  2129 => (x"48",x"00",x"00",x"08"),
  2130 => (x"74",x"54",x"54",x"5c"),
  2131 => (x"04",x"00",x"00",x"20"),
  2132 => (x"44",x"44",x"7f",x"3f"),
  2133 => (x"3c",x"00",x"00",x"00"),
  2134 => (x"7c",x"40",x"40",x"7c"),
  2135 => (x"1c",x"00",x"00",x"7c"),
  2136 => (x"3c",x"60",x"60",x"3c"),
  2137 => (x"7c",x"3c",x"00",x"1c"),
  2138 => (x"7c",x"60",x"30",x"60"),
  2139 => (x"6c",x"44",x"00",x"3c"),
  2140 => (x"6c",x"38",x"10",x"38"),
  2141 => (x"1c",x"00",x"00",x"44"),
  2142 => (x"3c",x"60",x"e0",x"bc"),
  2143 => (x"44",x"00",x"00",x"1c"),
  2144 => (x"4c",x"5c",x"74",x"64"),
  2145 => (x"08",x"00",x"00",x"44"),
  2146 => (x"41",x"77",x"3e",x"08"),
  2147 => (x"00",x"00",x"00",x"41"),
  2148 => (x"00",x"7f",x"7f",x"00"),
  2149 => (x"41",x"00",x"00",x"00"),
  2150 => (x"08",x"3e",x"77",x"41"),
  2151 => (x"01",x"02",x"00",x"08"),
  2152 => (x"02",x"02",x"03",x"01"),
  2153 => (x"7f",x"7f",x"00",x"01"),
  2154 => (x"7f",x"7f",x"7f",x"7f"),
  2155 => (x"08",x"08",x"00",x"7f"),
  2156 => (x"3e",x"3e",x"1c",x"1c"),
  2157 => (x"7f",x"7f",x"7f",x"7f"),
  2158 => (x"1c",x"1c",x"3e",x"3e"),
  2159 => (x"10",x"00",x"08",x"08"),
  2160 => (x"18",x"7c",x"7c",x"18"),
  2161 => (x"10",x"00",x"00",x"10"),
  2162 => (x"30",x"7c",x"7c",x"30"),
  2163 => (x"30",x"10",x"00",x"10"),
  2164 => (x"1e",x"78",x"60",x"60"),
  2165 => (x"66",x"42",x"00",x"06"),
  2166 => (x"66",x"3c",x"18",x"3c"),
  2167 => (x"38",x"78",x"00",x"42"),
  2168 => (x"6c",x"c6",x"c2",x"6a"),
  2169 => (x"00",x"60",x"00",x"38"),
  2170 => (x"00",x"00",x"60",x"00"),
  2171 => (x"5e",x"0e",x"00",x"60"),
  2172 => (x"0e",x"5d",x"5c",x"5b"),
  2173 => (x"c2",x"4c",x"71",x"1e"),
  2174 => (x"4b",x"bf",x"f6",x"eb"),
  2175 => (x"48",x"fa",x"eb",x"c2"),
  2176 => (x"f6",x"27",x"78",x"c0"),
  2177 => (x"bf",x"00",x"00",x"2a"),
  2178 => (x"99",x"49",x"bf",x"97"),
  2179 => (x"87",x"c8",x"c1",x"02"),
  2180 => (x"eb",x"c2",x"1e",x"c0"),
  2181 => (x"74",x"4d",x"bf",x"fa"),
  2182 => (x"87",x"c7",x"02",x"ad"),
  2183 => (x"c0",x"48",x"a6",x"c4"),
  2184 => (x"c4",x"87",x"c5",x"78"),
  2185 => (x"78",x"c1",x"48",x"a6"),
  2186 => (x"75",x"1e",x"66",x"c4"),
  2187 => (x"87",x"c4",x"ed",x"49"),
  2188 => (x"e0",x"c0",x"86",x"c8"),
  2189 => (x"87",x"f5",x"ee",x"49"),
  2190 => (x"6a",x"4a",x"a3",x"c4"),
  2191 => (x"87",x"f7",x"ef",x"49"),
  2192 => (x"c2",x"87",x"cd",x"f0"),
  2193 => (x"48",x"bf",x"fa",x"eb"),
  2194 => (x"eb",x"c2",x"80",x"c1"),
  2195 => (x"83",x"cc",x"58",x"fe"),
  2196 => (x"99",x"49",x"6b",x"97"),
  2197 => (x"87",x"f8",x"fe",x"05"),
  2198 => (x"bf",x"fa",x"eb",x"c2"),
  2199 => (x"ad",x"b7",x"c8",x"4d"),
  2200 => (x"c0",x"87",x"d9",x"03"),
  2201 => (x"eb",x"c2",x"1e",x"1e"),
  2202 => (x"ec",x"49",x"bf",x"fa"),
  2203 => (x"86",x"c8",x"87",x"c6"),
  2204 => (x"c1",x"87",x"dd",x"ef"),
  2205 => (x"ad",x"b7",x"c8",x"85"),
  2206 => (x"87",x"e7",x"ff",x"04"),
  2207 => (x"26",x"4d",x"26",x"26"),
  2208 => (x"26",x"4b",x"26",x"4c"),
  2209 => (x"4a",x"71",x"1e",x"4f"),
  2210 => (x"5a",x"fa",x"eb",x"c2"),
  2211 => (x"bf",x"fe",x"eb",x"c2"),
  2212 => (x"87",x"da",x"fd",x"49"),
  2213 => (x"bf",x"fa",x"eb",x"c2"),
  2214 => (x"c2",x"89",x"c1",x"49"),
  2215 => (x"71",x"59",x"c2",x"ec"),
  2216 => (x"26",x"87",x"cb",x"fd"),
  2217 => (x"c0",x"c1",x"1e",x"4f"),
  2218 => (x"87",x"d8",x"ea",x"49"),
  2219 => (x"48",x"eb",x"d6",x"c2"),
  2220 => (x"4f",x"26",x"78",x"c0"),
  2221 => (x"5c",x"5b",x"5e",x"0e"),
  2222 => (x"86",x"f4",x"0e",x"5d"),
  2223 => (x"c0",x"48",x"a6",x"c8"),
  2224 => (x"7e",x"bf",x"ec",x"78"),
  2225 => (x"eb",x"c2",x"80",x"fc"),
  2226 => (x"c2",x"78",x"bf",x"f6"),
  2227 => (x"4d",x"bf",x"c2",x"ec"),
  2228 => (x"c7",x"4c",x"bf",x"e8"),
  2229 => (x"87",x"f7",x"e5",x"49"),
  2230 => (x"99",x"c2",x"49",x"70"),
  2231 => (x"c2",x"87",x"cf",x"05"),
  2232 => (x"49",x"bf",x"e3",x"d6"),
  2233 => (x"99",x"6e",x"b9",x"ff"),
  2234 => (x"c0",x"02",x"99",x"c1"),
  2235 => (x"49",x"c7",x"87",x"ee"),
  2236 => (x"70",x"87",x"dc",x"e5"),
  2237 => (x"87",x"cd",x"02",x"98"),
  2238 => (x"c7",x"87",x"ca",x"e1"),
  2239 => (x"87",x"cf",x"e5",x"49"),
  2240 => (x"f3",x"05",x"98",x"70"),
  2241 => (x"eb",x"d6",x"c2",x"87"),
  2242 => (x"ba",x"c1",x"4a",x"bf"),
  2243 => (x"5a",x"ef",x"d6",x"c2"),
  2244 => (x"49",x"a2",x"c0",x"c1"),
  2245 => (x"c8",x"87",x"ed",x"e8"),
  2246 => (x"78",x"c1",x"48",x"a6"),
  2247 => (x"48",x"e3",x"d6",x"c2"),
  2248 => (x"d6",x"c2",x"78",x"6e"),
  2249 => (x"c1",x"05",x"bf",x"eb"),
  2250 => (x"a6",x"c4",x"87",x"da"),
  2251 => (x"c0",x"c0",x"c8",x"48"),
  2252 => (x"ef",x"d6",x"c2",x"78"),
  2253 => (x"bf",x"97",x"6e",x"7e"),
  2254 => (x"c1",x"48",x"6e",x"49"),
  2255 => (x"58",x"a6",x"c4",x"80"),
  2256 => (x"87",x"cb",x"e4",x"71"),
  2257 => (x"c3",x"02",x"98",x"70"),
  2258 => (x"b4",x"66",x"c4",x"87"),
  2259 => (x"c1",x"48",x"66",x"c4"),
  2260 => (x"a6",x"c8",x"28",x"b7"),
  2261 => (x"05",x"98",x"70",x"58"),
  2262 => (x"74",x"87",x"da",x"ff"),
  2263 => (x"99",x"ff",x"c3",x"49"),
  2264 => (x"49",x"c0",x"1e",x"71"),
  2265 => (x"74",x"87",x"d0",x"e6"),
  2266 => (x"29",x"b7",x"c8",x"49"),
  2267 => (x"49",x"c1",x"1e",x"71"),
  2268 => (x"c8",x"87",x"c4",x"e6"),
  2269 => (x"49",x"fd",x"c3",x"86"),
  2270 => (x"c3",x"87",x"d4",x"e3"),
  2271 => (x"ce",x"e3",x"49",x"fa"),
  2272 => (x"87",x"ca",x"c8",x"87"),
  2273 => (x"ff",x"c3",x"49",x"74"),
  2274 => (x"2c",x"b7",x"c8",x"99"),
  2275 => (x"9c",x"74",x"b4",x"71"),
  2276 => (x"ff",x"87",x"dd",x"02"),
  2277 => (x"6e",x"7e",x"bf",x"c8"),
  2278 => (x"e7",x"d6",x"c2",x"49"),
  2279 => (x"c0",x"c2",x"89",x"bf"),
  2280 => (x"87",x"c4",x"03",x"a9"),
  2281 => (x"87",x"ce",x"4c",x"c0"),
  2282 => (x"48",x"e7",x"d6",x"c2"),
  2283 => (x"87",x"c6",x"78",x"6e"),
  2284 => (x"48",x"e7",x"d6",x"c2"),
  2285 => (x"49",x"74",x"78",x"c0"),
  2286 => (x"ce",x"05",x"99",x"c8"),
  2287 => (x"49",x"f5",x"c3",x"87"),
  2288 => (x"70",x"87",x"cc",x"e2"),
  2289 => (x"02",x"99",x"c2",x"49"),
  2290 => (x"c2",x"87",x"ed",x"c0"),
  2291 => (x"02",x"bf",x"fe",x"eb"),
  2292 => (x"c1",x"48",x"87",x"c9"),
  2293 => (x"c2",x"ec",x"c2",x"88"),
  2294 => (x"c2",x"87",x"d8",x"58"),
  2295 => (x"49",x"bf",x"fa",x"eb"),
  2296 => (x"66",x"c4",x"91",x"cc"),
  2297 => (x"7e",x"a1",x"c8",x"81"),
  2298 => (x"c0",x"02",x"bf",x"6e"),
  2299 => (x"ff",x"4b",x"87",x"c5"),
  2300 => (x"c8",x"0f",x"73",x"49"),
  2301 => (x"78",x"c1",x"48",x"a6"),
  2302 => (x"99",x"c4",x"49",x"74"),
  2303 => (x"c3",x"87",x"ce",x"05"),
  2304 => (x"ca",x"e1",x"49",x"f2"),
  2305 => (x"c2",x"49",x"70",x"87"),
  2306 => (x"fd",x"c0",x"02",x"99"),
  2307 => (x"48",x"a6",x"c8",x"87"),
  2308 => (x"bf",x"fa",x"eb",x"c2"),
  2309 => (x"49",x"66",x"c8",x"78"),
  2310 => (x"eb",x"c2",x"89",x"c1"),
  2311 => (x"6e",x"7e",x"bf",x"fe"),
  2312 => (x"c0",x"06",x"a9",x"b7"),
  2313 => (x"c1",x"48",x"87",x"c9"),
  2314 => (x"c2",x"ec",x"c2",x"80"),
  2315 => (x"c8",x"87",x"d6",x"58"),
  2316 => (x"91",x"cc",x"49",x"66"),
  2317 => (x"c8",x"81",x"66",x"c4"),
  2318 => (x"bf",x"6e",x"7e",x"a1"),
  2319 => (x"87",x"c5",x"c0",x"02"),
  2320 => (x"73",x"49",x"fe",x"4b"),
  2321 => (x"48",x"a6",x"c8",x"0f"),
  2322 => (x"fd",x"c3",x"78",x"c1"),
  2323 => (x"fe",x"df",x"ff",x"49"),
  2324 => (x"c2",x"49",x"70",x"87"),
  2325 => (x"ee",x"c0",x"02",x"99"),
  2326 => (x"fe",x"eb",x"c2",x"87"),
  2327 => (x"c9",x"c0",x"02",x"bf"),
  2328 => (x"fe",x"eb",x"c2",x"87"),
  2329 => (x"c0",x"78",x"c0",x"48"),
  2330 => (x"eb",x"c2",x"87",x"d8"),
  2331 => (x"cc",x"49",x"bf",x"fa"),
  2332 => (x"81",x"66",x"c4",x"91"),
  2333 => (x"6e",x"7e",x"a1",x"c8"),
  2334 => (x"c5",x"c0",x"02",x"bf"),
  2335 => (x"49",x"fd",x"4b",x"87"),
  2336 => (x"a6",x"c8",x"0f",x"73"),
  2337 => (x"c3",x"78",x"c1",x"48"),
  2338 => (x"df",x"ff",x"49",x"fa"),
  2339 => (x"49",x"70",x"87",x"c1"),
  2340 => (x"c1",x"02",x"99",x"c2"),
  2341 => (x"a6",x"c8",x"87",x"c0"),
  2342 => (x"fa",x"eb",x"c2",x"48"),
  2343 => (x"66",x"c8",x"78",x"bf"),
  2344 => (x"c4",x"88",x"c1",x"48"),
  2345 => (x"eb",x"c2",x"58",x"a6"),
  2346 => (x"6e",x"48",x"bf",x"fe"),
  2347 => (x"c0",x"03",x"a8",x"b7"),
  2348 => (x"eb",x"c2",x"87",x"c9"),
  2349 => (x"78",x"6e",x"48",x"fe"),
  2350 => (x"c8",x"87",x"d6",x"c0"),
  2351 => (x"91",x"cc",x"49",x"66"),
  2352 => (x"c8",x"81",x"66",x"c4"),
  2353 => (x"bf",x"6e",x"7e",x"a1"),
  2354 => (x"87",x"c5",x"c0",x"02"),
  2355 => (x"73",x"49",x"fc",x"4b"),
  2356 => (x"48",x"a6",x"c8",x"0f"),
  2357 => (x"eb",x"c2",x"78",x"c1"),
  2358 => (x"c0",x"4a",x"bf",x"fe"),
  2359 => (x"c0",x"06",x"aa",x"b7"),
  2360 => (x"8a",x"c1",x"87",x"c9"),
  2361 => (x"01",x"aa",x"b7",x"c0"),
  2362 => (x"74",x"87",x"f7",x"ff"),
  2363 => (x"99",x"f0",x"c3",x"49"),
  2364 => (x"87",x"cf",x"c0",x"05"),
  2365 => (x"ff",x"49",x"da",x"c1"),
  2366 => (x"70",x"87",x"d4",x"dd"),
  2367 => (x"02",x"99",x"c2",x"49"),
  2368 => (x"c2",x"87",x"ce",x"c1"),
  2369 => (x"7e",x"bf",x"f6",x"eb"),
  2370 => (x"c2",x"48",x"a6",x"c4"),
  2371 => (x"78",x"bf",x"fe",x"eb"),
  2372 => (x"48",x"4a",x"66",x"c4"),
  2373 => (x"06",x"a8",x"b7",x"c0"),
  2374 => (x"6e",x"87",x"d0",x"c0"),
  2375 => (x"c4",x"80",x"cc",x"48"),
  2376 => (x"8a",x"c1",x"58",x"a6"),
  2377 => (x"01",x"aa",x"b7",x"c0"),
  2378 => (x"6e",x"87",x"f0",x"ff"),
  2379 => (x"c2",x"4b",x"bf",x"97"),
  2380 => (x"d1",x"c0",x"02",x"8b"),
  2381 => (x"c0",x"05",x"8b",x"87"),
  2382 => (x"4a",x"6e",x"87",x"d7"),
  2383 => (x"49",x"6a",x"82",x"c8"),
  2384 => (x"c0",x"87",x"c2",x"f5"),
  2385 => (x"4b",x"6e",x"87",x"cb"),
  2386 => (x"4b",x"6b",x"83",x"c8"),
  2387 => (x"73",x"49",x"66",x"c4"),
  2388 => (x"02",x"9d",x"75",x"0f"),
  2389 => (x"6d",x"87",x"e9",x"c0"),
  2390 => (x"87",x"e4",x"c0",x"02"),
  2391 => (x"db",x"ff",x"49",x"6d"),
  2392 => (x"49",x"70",x"87",x"ed"),
  2393 => (x"c0",x"02",x"99",x"c1"),
  2394 => (x"a5",x"c4",x"87",x"cb"),
  2395 => (x"fe",x"eb",x"c2",x"4b"),
  2396 => (x"4b",x"6b",x"49",x"bf"),
  2397 => (x"02",x"85",x"c8",x"0f"),
  2398 => (x"6d",x"87",x"c5",x"c0"),
  2399 => (x"87",x"dc",x"ff",x"05"),
  2400 => (x"c0",x"02",x"66",x"c8"),
  2401 => (x"eb",x"c2",x"87",x"c8"),
  2402 => (x"f1",x"49",x"bf",x"fe"),
  2403 => (x"8e",x"f4",x"87",x"e0"),
  2404 => (x"58",x"87",x"ea",x"f3"),
  2405 => (x"1d",x"14",x"11",x"12"),
  2406 => (x"5a",x"23",x"1c",x"1b"),
  2407 => (x"f5",x"94",x"91",x"59"),
  2408 => (x"00",x"f4",x"eb",x"f2"),
  2409 => (x"00",x"00",x"00",x"00"),
  2410 => (x"00",x"00",x"00",x"00"),
  2411 => (x"58",x"00",x"00",x"00"),
  2412 => (x"1d",x"11",x"14",x"12"),
  2413 => (x"5a",x"23",x"1c",x"1b"),
  2414 => (x"f5",x"91",x"94",x"59"),
  2415 => (x"00",x"f4",x"eb",x"f2"),
  2416 => (x"00",x"00",x"25",x"c4"),
  2417 => (x"4f",x"54",x"55",x"41"),
  2418 => (x"54",x"4f",x"4f",x"42"),
  2419 => (x"00",x"53",x"45",x"4e"),
  2420 => (x"00",x"00",x"19",x"c4"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

