
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"e7",x"c2",x"87"),
    12 => (x"48",x"c0",x"c4",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"05",x"88"),
    17 => (x"49",x"dc",x"e7",x"c2"),
    18 => (x"48",x"ec",x"d2",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"ea",x"d2",x"c2",x"87"),
    25 => (x"e6",x"d2",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e0",x"c1",x"87",x"f7"),
    29 => (x"d2",x"c2",x"87",x"d9"),
    30 => (x"d2",x"c2",x"4d",x"ea"),
    31 => (x"ad",x"74",x"4c",x"ea"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"c0",x"4b",x"71",x"0e"),
    37 => (x"9a",x"4a",x"13",x"4c"),
    38 => (x"72",x"87",x"cd",x"02"),
    39 => (x"87",x"e0",x"c0",x"49"),
    40 => (x"4a",x"13",x"84",x"c1"),
    41 => (x"87",x"f3",x"05",x"9a"),
    42 => (x"4c",x"26",x"48",x"74"),
    43 => (x"4f",x"26",x"4b",x"26"),
    44 => (x"81",x"48",x"73",x"1e"),
    45 => (x"c5",x"02",x"a9",x"73"),
    46 => (x"05",x"53",x"12",x"87"),
    47 => (x"4f",x"26",x"87",x"f6"),
    48 => (x"c0",x"ff",x"1e",x"1e"),
    49 => (x"c4",x"48",x"6a",x"4a"),
    50 => (x"a6",x"c4",x"98",x"c0"),
    51 => (x"02",x"98",x"70",x"58"),
    52 => (x"7a",x"71",x"87",x"f3"),
    53 => (x"4f",x"26",x"26",x"48"),
    54 => (x"ff",x"1e",x"73",x"1e"),
    55 => (x"ff",x"c3",x"4b",x"d4"),
    56 => (x"c3",x"4a",x"6b",x"7b"),
    57 => (x"49",x"6b",x"7b",x"ff"),
    58 => (x"b1",x"72",x"32",x"c8"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"71",x"31",x"c8",x"4a"),
    61 => (x"7b",x"ff",x"c3",x"b2"),
    62 => (x"32",x"c8",x"49",x"6b"),
    63 => (x"48",x"71",x"b1",x"72"),
    64 => (x"4d",x"26",x"87",x"c4"),
    65 => (x"4b",x"26",x"4c",x"26"),
    66 => (x"5e",x"0e",x"4f",x"26"),
    67 => (x"0e",x"5d",x"5c",x"5b"),
    68 => (x"d4",x"ff",x"4a",x"71"),
    69 => (x"c3",x"48",x"72",x"4c"),
    70 => (x"7c",x"70",x"98",x"ff"),
    71 => (x"bf",x"ec",x"d2",x"c2"),
    72 => (x"d0",x"87",x"c8",x"05"),
    73 => (x"30",x"c9",x"48",x"66"),
    74 => (x"d0",x"58",x"a6",x"d4"),
    75 => (x"29",x"d8",x"49",x"66"),
    76 => (x"ff",x"c3",x"48",x"71"),
    77 => (x"d0",x"7c",x"70",x"98"),
    78 => (x"29",x"d0",x"49",x"66"),
    79 => (x"ff",x"c3",x"48",x"71"),
    80 => (x"d0",x"7c",x"70",x"98"),
    81 => (x"29",x"c8",x"49",x"66"),
    82 => (x"ff",x"c3",x"48",x"71"),
    83 => (x"d0",x"7c",x"70",x"98"),
    84 => (x"ff",x"c3",x"48",x"66"),
    85 => (x"72",x"7c",x"70",x"98"),
    86 => (x"71",x"29",x"d0",x"49"),
    87 => (x"98",x"ff",x"c3",x"48"),
    88 => (x"4b",x"6c",x"7c",x"70"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"ff",x"fd"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"df",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c1",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"de",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"49",x"e3",x"c8",x"78"),
   125 => (x"d3",x"87",x"d5",x"fa"),
   126 => (x"c0",x"1e",x"c0",x"4b"),
   127 => (x"c1",x"c1",x"f0",x"ff"),
   128 => (x"87",x"c6",x"fc",x"49"),
   129 => (x"98",x"70",x"86",x"c4"),
   130 => (x"ff",x"87",x"ca",x"05"),
   131 => (x"ff",x"c3",x"48",x"d4"),
   132 => (x"cb",x"48",x"c1",x"78"),
   133 => (x"87",x"eb",x"fd",x"87"),
   134 => (x"ff",x"05",x"8b",x"c1"),
   135 => (x"48",x"c0",x"87",x"db"),
   136 => (x"43",x"87",x"e3",x"fb"),
   137 => (x"53",x"00",x"44",x"4d"),
   138 => (x"20",x"43",x"48",x"44"),
   139 => (x"6c",x"69",x"61",x"66"),
   140 => (x"49",x"00",x"0a",x"21"),
   141 => (x"00",x"52",x"52",x"45"),
   142 => (x"00",x"49",x"50",x"53"),
   143 => (x"74",x"69",x"72",x"57"),
   144 => (x"61",x"66",x"20",x"65"),
   145 => (x"64",x"65",x"6c",x"69"),
   146 => (x"5e",x"0e",x"00",x"0a"),
   147 => (x"ff",x"0e",x"5c",x"5b"),
   148 => (x"ee",x"fc",x"4c",x"d4"),
   149 => (x"1e",x"ea",x"c6",x"87"),
   150 => (x"c1",x"f0",x"e1",x"c0"),
   151 => (x"e9",x"fa",x"49",x"c8"),
   152 => (x"c1",x"86",x"c4",x"87"),
   153 => (x"87",x"c8",x"02",x"a8"),
   154 => (x"c0",x"87",x"fd",x"fd"),
   155 => (x"87",x"e8",x"c1",x"48"),
   156 => (x"70",x"87",x"e5",x"f9"),
   157 => (x"ff",x"ff",x"cf",x"49"),
   158 => (x"a9",x"ea",x"c6",x"99"),
   159 => (x"fd",x"87",x"c8",x"02"),
   160 => (x"48",x"c0",x"87",x"e6"),
   161 => (x"c3",x"87",x"d1",x"c1"),
   162 => (x"f1",x"c0",x"7c",x"ff"),
   163 => (x"87",x"c7",x"fc",x"4b"),
   164 => (x"c0",x"02",x"98",x"70"),
   165 => (x"1e",x"c0",x"87",x"eb"),
   166 => (x"c1",x"f0",x"ff",x"c0"),
   167 => (x"e9",x"f9",x"49",x"fa"),
   168 => (x"70",x"86",x"c4",x"87"),
   169 => (x"87",x"d9",x"05",x"98"),
   170 => (x"6c",x"7c",x"ff",x"c3"),
   171 => (x"7c",x"ff",x"c3",x"49"),
   172 => (x"c1",x"7c",x"7c",x"7c"),
   173 => (x"c4",x"02",x"99",x"c0"),
   174 => (x"db",x"48",x"c1",x"87"),
   175 => (x"d7",x"48",x"c0",x"87"),
   176 => (x"05",x"ab",x"c2",x"87"),
   177 => (x"e7",x"c8",x"87",x"ca"),
   178 => (x"87",x"c0",x"f7",x"49"),
   179 => (x"87",x"c8",x"48",x"c0"),
   180 => (x"fe",x"05",x"8b",x"c1"),
   181 => (x"48",x"c0",x"87",x"f7"),
   182 => (x"0e",x"87",x"e9",x"f8"),
   183 => (x"5d",x"5c",x"5b",x"5e"),
   184 => (x"d0",x"ff",x"1e",x"0e"),
   185 => (x"c0",x"c0",x"c8",x"4d"),
   186 => (x"ec",x"d2",x"c2",x"4b"),
   187 => (x"c8",x"78",x"c1",x"48"),
   188 => (x"d7",x"f6",x"49",x"f8"),
   189 => (x"6d",x"4c",x"c7",x"87"),
   190 => (x"c4",x"98",x"73",x"48"),
   191 => (x"98",x"70",x"58",x"a6"),
   192 => (x"6d",x"87",x"cc",x"02"),
   193 => (x"c4",x"98",x"73",x"48"),
   194 => (x"98",x"70",x"58",x"a6"),
   195 => (x"c2",x"87",x"f4",x"05"),
   196 => (x"87",x"ef",x"f9",x"7d"),
   197 => (x"98",x"73",x"48",x"6d"),
   198 => (x"70",x"58",x"a6",x"c4"),
   199 => (x"87",x"cc",x"02",x"98"),
   200 => (x"98",x"73",x"48",x"6d"),
   201 => (x"70",x"58",x"a6",x"c4"),
   202 => (x"87",x"f4",x"05",x"98"),
   203 => (x"1e",x"c0",x"7d",x"c3"),
   204 => (x"c1",x"d0",x"e5",x"c0"),
   205 => (x"d1",x"f7",x"49",x"c0"),
   206 => (x"c1",x"86",x"c4",x"87"),
   207 => (x"87",x"c1",x"05",x"a8"),
   208 => (x"05",x"ac",x"c2",x"4c"),
   209 => (x"f3",x"c8",x"87",x"cb"),
   210 => (x"87",x"c0",x"f5",x"49"),
   211 => (x"ce",x"c1",x"48",x"c0"),
   212 => (x"05",x"8c",x"c1",x"87"),
   213 => (x"fb",x"87",x"e0",x"fe"),
   214 => (x"d2",x"c2",x"87",x"f0"),
   215 => (x"98",x"70",x"58",x"f0"),
   216 => (x"c1",x"87",x"cd",x"05"),
   217 => (x"f0",x"ff",x"c0",x"1e"),
   218 => (x"f6",x"49",x"d0",x"c1"),
   219 => (x"86",x"c4",x"87",x"dc"),
   220 => (x"c3",x"48",x"d4",x"ff"),
   221 => (x"dd",x"c5",x"78",x"ff"),
   222 => (x"f4",x"d2",x"c2",x"87"),
   223 => (x"73",x"48",x"6d",x"58"),
   224 => (x"58",x"a6",x"c4",x"98"),
   225 => (x"cc",x"02",x"98",x"70"),
   226 => (x"73",x"48",x"6d",x"87"),
   227 => (x"58",x"a6",x"c4",x"98"),
   228 => (x"f4",x"05",x"98",x"70"),
   229 => (x"ff",x"7d",x"c2",x"87"),
   230 => (x"ff",x"c3",x"48",x"d4"),
   231 => (x"26",x"48",x"c1",x"78"),
   232 => (x"0e",x"87",x"df",x"f5"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"c8",x"1e",x"0e"),
   235 => (x"4c",x"c0",x"4b",x"c0"),
   236 => (x"df",x"cd",x"ee",x"c5"),
   237 => (x"5c",x"a6",x"c4",x"4a"),
   238 => (x"c3",x"4c",x"d4",x"ff"),
   239 => (x"48",x"6c",x"7c",x"ff"),
   240 => (x"05",x"a8",x"fe",x"c3"),
   241 => (x"71",x"87",x"c0",x"c2"),
   242 => (x"e2",x"c0",x"05",x"99"),
   243 => (x"bf",x"d0",x"ff",x"87"),
   244 => (x"c4",x"98",x"73",x"48"),
   245 => (x"98",x"70",x"58",x"a6"),
   246 => (x"ff",x"87",x"ce",x"02"),
   247 => (x"73",x"48",x"bf",x"d0"),
   248 => (x"58",x"a6",x"c4",x"98"),
   249 => (x"f2",x"05",x"98",x"70"),
   250 => (x"48",x"d0",x"ff",x"87"),
   251 => (x"d4",x"78",x"d1",x"c4"),
   252 => (x"b7",x"c0",x"48",x"66"),
   253 => (x"e0",x"c0",x"06",x"a8"),
   254 => (x"7c",x"ff",x"c3",x"87"),
   255 => (x"99",x"71",x"4a",x"6c"),
   256 => (x"71",x"87",x"c7",x"02"),
   257 => (x"0a",x"7a",x"97",x"0a"),
   258 => (x"66",x"d4",x"81",x"c1"),
   259 => (x"d8",x"88",x"c1",x"48"),
   260 => (x"b7",x"c0",x"58",x"a6"),
   261 => (x"e0",x"ff",x"01",x"a8"),
   262 => (x"7c",x"ff",x"c3",x"87"),
   263 => (x"05",x"99",x"71",x"7c"),
   264 => (x"ff",x"87",x"e1",x"c0"),
   265 => (x"73",x"48",x"bf",x"d0"),
   266 => (x"58",x"a6",x"c4",x"98"),
   267 => (x"ce",x"02",x"98",x"70"),
   268 => (x"bf",x"d0",x"ff",x"87"),
   269 => (x"c4",x"98",x"73",x"48"),
   270 => (x"98",x"70",x"58",x"a6"),
   271 => (x"ff",x"87",x"f2",x"05"),
   272 => (x"78",x"d0",x"48",x"d0"),
   273 => (x"c1",x"7e",x"4a",x"c1"),
   274 => (x"ee",x"fd",x"05",x"8a"),
   275 => (x"26",x"48",x"6e",x"87"),
   276 => (x"0e",x"87",x"ef",x"f2"),
   277 => (x"0e",x"5c",x"5b",x"5e"),
   278 => (x"c8",x"4a",x"71",x"1e"),
   279 => (x"c0",x"4b",x"c0",x"c0"),
   280 => (x"48",x"d4",x"ff",x"4c"),
   281 => (x"ff",x"78",x"ff",x"c3"),
   282 => (x"73",x"48",x"bf",x"d0"),
   283 => (x"58",x"a6",x"c4",x"98"),
   284 => (x"ce",x"02",x"98",x"70"),
   285 => (x"bf",x"d0",x"ff",x"87"),
   286 => (x"c4",x"98",x"73",x"48"),
   287 => (x"98",x"70",x"58",x"a6"),
   288 => (x"ff",x"87",x"f2",x"05"),
   289 => (x"c3",x"c4",x"48",x"d0"),
   290 => (x"48",x"d4",x"ff",x"78"),
   291 => (x"72",x"78",x"ff",x"c3"),
   292 => (x"f0",x"ff",x"c0",x"1e"),
   293 => (x"f1",x"49",x"d1",x"c1"),
   294 => (x"86",x"c4",x"87",x"f0"),
   295 => (x"c0",x"05",x"98",x"70"),
   296 => (x"c0",x"c8",x"87",x"ee"),
   297 => (x"49",x"66",x"d4",x"1e"),
   298 => (x"c4",x"87",x"f8",x"fb"),
   299 => (x"ff",x"4c",x"70",x"86"),
   300 => (x"73",x"48",x"bf",x"d0"),
   301 => (x"58",x"a6",x"c4",x"98"),
   302 => (x"ce",x"02",x"98",x"70"),
   303 => (x"bf",x"d0",x"ff",x"87"),
   304 => (x"c4",x"98",x"73",x"48"),
   305 => (x"98",x"70",x"58",x"a6"),
   306 => (x"ff",x"87",x"f2",x"05"),
   307 => (x"78",x"c2",x"48",x"d0"),
   308 => (x"f0",x"26",x"48",x"74"),
   309 => (x"5e",x"0e",x"87",x"ee"),
   310 => (x"0e",x"5d",x"5c",x"5b"),
   311 => (x"ff",x"c0",x"1e",x"c0"),
   312 => (x"49",x"c9",x"c1",x"f0"),
   313 => (x"d2",x"87",x"e3",x"f0"),
   314 => (x"fa",x"d2",x"c2",x"1e"),
   315 => (x"87",x"f3",x"fa",x"49"),
   316 => (x"4c",x"c0",x"86",x"c8"),
   317 => (x"b7",x"d2",x"84",x"c1"),
   318 => (x"87",x"f8",x"04",x"ac"),
   319 => (x"97",x"fa",x"d2",x"c2"),
   320 => (x"c0",x"c3",x"49",x"bf"),
   321 => (x"a9",x"c0",x"c1",x"99"),
   322 => (x"87",x"e7",x"c0",x"05"),
   323 => (x"97",x"c1",x"d3",x"c2"),
   324 => (x"31",x"d0",x"49",x"bf"),
   325 => (x"97",x"c2",x"d3",x"c2"),
   326 => (x"32",x"c8",x"4a",x"bf"),
   327 => (x"d3",x"c2",x"b1",x"72"),
   328 => (x"4a",x"bf",x"97",x"c3"),
   329 => (x"cf",x"4c",x"71",x"b1"),
   330 => (x"9c",x"ff",x"ff",x"ff"),
   331 => (x"34",x"ca",x"84",x"c1"),
   332 => (x"c2",x"87",x"e7",x"c1"),
   333 => (x"bf",x"97",x"c3",x"d3"),
   334 => (x"c6",x"31",x"c1",x"49"),
   335 => (x"c4",x"d3",x"c2",x"99"),
   336 => (x"c7",x"4a",x"bf",x"97"),
   337 => (x"b1",x"72",x"2a",x"b7"),
   338 => (x"97",x"ff",x"d2",x"c2"),
   339 => (x"cf",x"4d",x"4a",x"bf"),
   340 => (x"c0",x"d3",x"c2",x"9d"),
   341 => (x"c3",x"4a",x"bf",x"97"),
   342 => (x"c2",x"32",x"ca",x"9a"),
   343 => (x"bf",x"97",x"c1",x"d3"),
   344 => (x"73",x"33",x"c2",x"4b"),
   345 => (x"c2",x"d3",x"c2",x"b2"),
   346 => (x"c3",x"4b",x"bf",x"97"),
   347 => (x"b7",x"c6",x"9b",x"c0"),
   348 => (x"c2",x"b2",x"73",x"2b"),
   349 => (x"71",x"48",x"c1",x"81"),
   350 => (x"c1",x"49",x"70",x"30"),
   351 => (x"70",x"30",x"75",x"48"),
   352 => (x"c1",x"4c",x"72",x"4d"),
   353 => (x"c8",x"94",x"71",x"84"),
   354 => (x"06",x"ad",x"b7",x"c0"),
   355 => (x"34",x"c1",x"87",x"cc"),
   356 => (x"c0",x"c8",x"2d",x"b7"),
   357 => (x"ff",x"01",x"ad",x"b7"),
   358 => (x"48",x"74",x"87",x"f4"),
   359 => (x"0e",x"87",x"e3",x"ed"),
   360 => (x"0e",x"5c",x"5b",x"5e"),
   361 => (x"4c",x"c0",x"4b",x"71"),
   362 => (x"c0",x"48",x"66",x"d0"),
   363 => (x"c0",x"06",x"a8",x"b7"),
   364 => (x"4a",x"13",x"87",x"e3"),
   365 => (x"bf",x"97",x"66",x"cc"),
   366 => (x"48",x"66",x"cc",x"49"),
   367 => (x"a6",x"d0",x"80",x"c1"),
   368 => (x"aa",x"b7",x"71",x"58"),
   369 => (x"c1",x"87",x"c4",x"02"),
   370 => (x"c1",x"87",x"cc",x"48"),
   371 => (x"b7",x"66",x"d0",x"84"),
   372 => (x"dd",x"ff",x"04",x"ac"),
   373 => (x"c2",x"48",x"c0",x"87"),
   374 => (x"26",x"4d",x"26",x"87"),
   375 => (x"26",x"4b",x"26",x"4c"),
   376 => (x"5b",x"5e",x"0e",x"4f"),
   377 => (x"c2",x"0e",x"5d",x"5c"),
   378 => (x"c0",x"48",x"e0",x"db"),
   379 => (x"d8",x"d3",x"c2",x"78"),
   380 => (x"f9",x"49",x"c0",x"1e"),
   381 => (x"86",x"c4",x"87",x"dd"),
   382 => (x"c5",x"05",x"98",x"70"),
   383 => (x"c8",x"48",x"c0",x"87"),
   384 => (x"4b",x"c0",x"87",x"ef"),
   385 => (x"48",x"d8",x"e0",x"c2"),
   386 => (x"1e",x"c8",x"78",x"c1"),
   387 => (x"1e",x"fd",x"e0",x"c0"),
   388 => (x"49",x"ce",x"d4",x"c2"),
   389 => (x"c8",x"87",x"c8",x"fe"),
   390 => (x"05",x"98",x"70",x"86"),
   391 => (x"e0",x"c2",x"87",x"c6"),
   392 => (x"78",x"c0",x"48",x"d8"),
   393 => (x"e1",x"c0",x"1e",x"c8"),
   394 => (x"d4",x"c2",x"1e",x"c6"),
   395 => (x"ee",x"fd",x"49",x"ea"),
   396 => (x"70",x"86",x"c8",x"87"),
   397 => (x"87",x"c6",x"05",x"98"),
   398 => (x"48",x"d8",x"e0",x"c2"),
   399 => (x"e0",x"c2",x"78",x"c0"),
   400 => (x"c0",x"02",x"bf",x"d8"),
   401 => (x"da",x"c2",x"87",x"fa"),
   402 => (x"c2",x"4b",x"bf",x"de"),
   403 => (x"bf",x"9f",x"d6",x"db"),
   404 => (x"ea",x"d6",x"c5",x"4a"),
   405 => (x"87",x"c7",x"05",x"aa"),
   406 => (x"bf",x"de",x"da",x"c2"),
   407 => (x"ca",x"87",x"cc",x"4b"),
   408 => (x"02",x"aa",x"d5",x"e9"),
   409 => (x"48",x"c0",x"87",x"c5"),
   410 => (x"c2",x"87",x"c6",x"c7"),
   411 => (x"73",x"1e",x"d8",x"d3"),
   412 => (x"87",x"df",x"f7",x"49"),
   413 => (x"98",x"70",x"86",x"c4"),
   414 => (x"c0",x"87",x"c5",x"05"),
   415 => (x"87",x"f1",x"c6",x"48"),
   416 => (x"e1",x"c0",x"1e",x"c8"),
   417 => (x"d4",x"c2",x"1e",x"cf"),
   418 => (x"d2",x"fc",x"49",x"ea"),
   419 => (x"70",x"86",x"c8",x"87"),
   420 => (x"87",x"c8",x"05",x"98"),
   421 => (x"48",x"e0",x"db",x"c2"),
   422 => (x"87",x"da",x"78",x"c1"),
   423 => (x"e1",x"c0",x"1e",x"c8"),
   424 => (x"d4",x"c2",x"1e",x"d8"),
   425 => (x"f6",x"fb",x"49",x"ce"),
   426 => (x"70",x"86",x"c8",x"87"),
   427 => (x"c5",x"c0",x"02",x"98"),
   428 => (x"c5",x"48",x"c0",x"87"),
   429 => (x"db",x"c2",x"87",x"fb"),
   430 => (x"49",x"bf",x"97",x"d6"),
   431 => (x"05",x"a9",x"d5",x"c1"),
   432 => (x"c2",x"87",x"cd",x"c0"),
   433 => (x"bf",x"97",x"d7",x"db"),
   434 => (x"a9",x"ea",x"c2",x"49"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dc",x"c5",x"48",x"c0"),
   437 => (x"d8",x"d3",x"c2",x"87"),
   438 => (x"c3",x"4c",x"bf",x"97"),
   439 => (x"c0",x"02",x"ac",x"e9"),
   440 => (x"eb",x"c3",x"87",x"cc"),
   441 => (x"c5",x"c0",x"02",x"ac"),
   442 => (x"c5",x"48",x"c0",x"87"),
   443 => (x"d3",x"c2",x"87",x"c3"),
   444 => (x"49",x"bf",x"97",x"e3"),
   445 => (x"cc",x"c0",x"05",x"99"),
   446 => (x"e4",x"d3",x"c2",x"87"),
   447 => (x"c2",x"49",x"bf",x"97"),
   448 => (x"c5",x"c0",x"02",x"a9"),
   449 => (x"c4",x"48",x"c0",x"87"),
   450 => (x"d3",x"c2",x"87",x"e7"),
   451 => (x"48",x"bf",x"97",x"e5"),
   452 => (x"58",x"dc",x"db",x"c2"),
   453 => (x"db",x"c2",x"88",x"c1"),
   454 => (x"d3",x"c2",x"58",x"e0"),
   455 => (x"49",x"bf",x"97",x"e6"),
   456 => (x"d3",x"c2",x"81",x"73"),
   457 => (x"4a",x"bf",x"97",x"e7"),
   458 => (x"71",x"35",x"c8",x"4d"),
   459 => (x"f8",x"df",x"c2",x"85"),
   460 => (x"e8",x"d3",x"c2",x"5d"),
   461 => (x"c2",x"48",x"bf",x"97"),
   462 => (x"c2",x"58",x"cc",x"e0"),
   463 => (x"02",x"bf",x"e0",x"db"),
   464 => (x"c8",x"87",x"dc",x"c2"),
   465 => (x"f4",x"e0",x"c0",x"1e"),
   466 => (x"ea",x"d4",x"c2",x"1e"),
   467 => (x"87",x"cf",x"f9",x"49"),
   468 => (x"98",x"70",x"86",x"c8"),
   469 => (x"87",x"c5",x"c0",x"02"),
   470 => (x"d4",x"c3",x"48",x"c0"),
   471 => (x"d8",x"db",x"c2",x"87"),
   472 => (x"c4",x"48",x"4a",x"bf"),
   473 => (x"e8",x"db",x"c2",x"30"),
   474 => (x"c8",x"e0",x"c2",x"58"),
   475 => (x"fd",x"d3",x"c2",x"5a"),
   476 => (x"c8",x"49",x"bf",x"97"),
   477 => (x"fc",x"d3",x"c2",x"31"),
   478 => (x"a1",x"4b",x"bf",x"97"),
   479 => (x"fe",x"d3",x"c2",x"49"),
   480 => (x"d0",x"4b",x"bf",x"97"),
   481 => (x"49",x"a1",x"73",x"33"),
   482 => (x"97",x"ff",x"d3",x"c2"),
   483 => (x"33",x"d8",x"4b",x"bf"),
   484 => (x"c2",x"49",x"a1",x"73"),
   485 => (x"c2",x"59",x"d0",x"e0"),
   486 => (x"91",x"bf",x"c8",x"e0"),
   487 => (x"bf",x"f4",x"df",x"c2"),
   488 => (x"fc",x"df",x"c2",x"81"),
   489 => (x"c5",x"d4",x"c2",x"59"),
   490 => (x"c8",x"4b",x"bf",x"97"),
   491 => (x"c4",x"d4",x"c2",x"33"),
   492 => (x"a3",x"4c",x"bf",x"97"),
   493 => (x"c6",x"d4",x"c2",x"4b"),
   494 => (x"d0",x"4c",x"bf",x"97"),
   495 => (x"4b",x"a3",x"74",x"34"),
   496 => (x"97",x"c7",x"d4",x"c2"),
   497 => (x"9c",x"cf",x"4c",x"bf"),
   498 => (x"a3",x"74",x"34",x"d8"),
   499 => (x"c0",x"e0",x"c2",x"4b"),
   500 => (x"73",x"8b",x"c2",x"5b"),
   501 => (x"c0",x"e0",x"c2",x"92"),
   502 => (x"78",x"a1",x"72",x"48"),
   503 => (x"c2",x"87",x"cb",x"c1"),
   504 => (x"bf",x"97",x"ea",x"d3"),
   505 => (x"c2",x"31",x"c8",x"49"),
   506 => (x"bf",x"97",x"e9",x"d3"),
   507 => (x"c2",x"49",x"a1",x"4a"),
   508 => (x"c5",x"59",x"e8",x"db"),
   509 => (x"81",x"ff",x"c7",x"31"),
   510 => (x"e0",x"c2",x"29",x"c9"),
   511 => (x"d3",x"c2",x"59",x"c8"),
   512 => (x"4a",x"bf",x"97",x"ef"),
   513 => (x"d3",x"c2",x"32",x"c8"),
   514 => (x"4b",x"bf",x"97",x"ee"),
   515 => (x"e0",x"c2",x"4a",x"a2"),
   516 => (x"e0",x"c2",x"5a",x"d0"),
   517 => (x"75",x"92",x"bf",x"c8"),
   518 => (x"c4",x"e0",x"c2",x"82"),
   519 => (x"fc",x"df",x"c2",x"5a"),
   520 => (x"c2",x"78",x"c0",x"48"),
   521 => (x"72",x"48",x"f8",x"df"),
   522 => (x"49",x"c0",x"78",x"a1"),
   523 => (x"c1",x"87",x"f7",x"c7"),
   524 => (x"87",x"e5",x"f6",x"48"),
   525 => (x"33",x"54",x"41",x"46"),
   526 => (x"20",x"20",x"20",x"32"),
   527 => (x"54",x"41",x"46",x"00"),
   528 => (x"20",x"20",x"36",x"31"),
   529 => (x"41",x"46",x"00",x"20"),
   530 => (x"20",x"32",x"33",x"54"),
   531 => (x"46",x"00",x"20",x"20"),
   532 => (x"32",x"33",x"54",x"41"),
   533 => (x"00",x"20",x"20",x"20"),
   534 => (x"31",x"54",x"41",x"46"),
   535 => (x"20",x"20",x"20",x"36"),
   536 => (x"5b",x"5e",x"0e",x"00"),
   537 => (x"71",x"0e",x"5d",x"5c"),
   538 => (x"e0",x"db",x"c2",x"4a"),
   539 => (x"87",x"cc",x"02",x"bf"),
   540 => (x"b7",x"c7",x"4b",x"72"),
   541 => (x"c1",x"4d",x"72",x"2b"),
   542 => (x"87",x"ca",x"9d",x"ff"),
   543 => (x"b7",x"c8",x"4b",x"72"),
   544 => (x"c3",x"4d",x"72",x"2b"),
   545 => (x"d3",x"c2",x"9d",x"ff"),
   546 => (x"df",x"c2",x"1e",x"d8"),
   547 => (x"73",x"49",x"bf",x"f4"),
   548 => (x"fe",x"ee",x"71",x"81"),
   549 => (x"70",x"86",x"c4",x"87"),
   550 => (x"87",x"c5",x"05",x"98"),
   551 => (x"e6",x"c0",x"48",x"c0"),
   552 => (x"e0",x"db",x"c2",x"87"),
   553 => (x"87",x"d2",x"02",x"bf"),
   554 => (x"91",x"c4",x"49",x"75"),
   555 => (x"81",x"d8",x"d3",x"c2"),
   556 => (x"ff",x"cf",x"4c",x"69"),
   557 => (x"9c",x"ff",x"ff",x"ff"),
   558 => (x"49",x"75",x"87",x"cb"),
   559 => (x"d3",x"c2",x"91",x"c2"),
   560 => (x"69",x"9f",x"81",x"d8"),
   561 => (x"f4",x"48",x"74",x"4c"),
   562 => (x"5e",x"0e",x"87",x"cf"),
   563 => (x"0e",x"5d",x"5c",x"5b"),
   564 => (x"4c",x"71",x"86",x"f4"),
   565 => (x"e0",x"c2",x"4b",x"c0"),
   566 => (x"c4",x"7e",x"bf",x"d0"),
   567 => (x"e0",x"c2",x"48",x"a6"),
   568 => (x"c8",x"78",x"bf",x"d4"),
   569 => (x"78",x"c0",x"48",x"a6"),
   570 => (x"bf",x"e4",x"db",x"c2"),
   571 => (x"06",x"a8",x"c0",x"48"),
   572 => (x"c8",x"87",x"dd",x"c2"),
   573 => (x"99",x"cf",x"49",x"66"),
   574 => (x"c2",x"87",x"d8",x"05"),
   575 => (x"c8",x"1e",x"d8",x"d3"),
   576 => (x"c1",x"48",x"49",x"66"),
   577 => (x"58",x"a6",x"cc",x"80"),
   578 => (x"c4",x"87",x"c8",x"ed"),
   579 => (x"d8",x"d3",x"c2",x"86"),
   580 => (x"c0",x"87",x"c3",x"4b"),
   581 => (x"6b",x"97",x"83",x"e0"),
   582 => (x"c1",x"02",x"9a",x"4a"),
   583 => (x"e5",x"c3",x"87",x"e1"),
   584 => (x"da",x"c1",x"02",x"aa"),
   585 => (x"49",x"a3",x"cb",x"87"),
   586 => (x"d8",x"49",x"69",x"97"),
   587 => (x"ce",x"c1",x"05",x"99"),
   588 => (x"c0",x"1e",x"cb",x"87"),
   589 => (x"73",x"1e",x"66",x"e0"),
   590 => (x"87",x"e3",x"f1",x"49"),
   591 => (x"98",x"70",x"86",x"c8"),
   592 => (x"87",x"fb",x"c0",x"05"),
   593 => (x"c4",x"4a",x"a3",x"dc"),
   594 => (x"79",x"6a",x"49",x"a4"),
   595 => (x"c8",x"49",x"a3",x"da"),
   596 => (x"69",x"9f",x"4d",x"a4"),
   597 => (x"db",x"c2",x"7d",x"48"),
   598 => (x"d3",x"02",x"bf",x"e0"),
   599 => (x"49",x"a3",x"d4",x"87"),
   600 => (x"c0",x"49",x"69",x"9f"),
   601 => (x"71",x"99",x"ff",x"ff"),
   602 => (x"c4",x"30",x"d0",x"48"),
   603 => (x"87",x"c2",x"58",x"a6"),
   604 => (x"48",x"6e",x"7e",x"c0"),
   605 => (x"7d",x"70",x"80",x"6d"),
   606 => (x"48",x"c1",x"7c",x"c0"),
   607 => (x"c8",x"87",x"c5",x"c1"),
   608 => (x"80",x"c1",x"48",x"66"),
   609 => (x"c2",x"58",x"a6",x"cc"),
   610 => (x"a8",x"bf",x"e4",x"db"),
   611 => (x"87",x"e3",x"fd",x"04"),
   612 => (x"bf",x"e0",x"db",x"c2"),
   613 => (x"87",x"ea",x"c0",x"02"),
   614 => (x"c4",x"fb",x"49",x"6e"),
   615 => (x"58",x"a6",x"c4",x"87"),
   616 => (x"ff",x"cf",x"49",x"70"),
   617 => (x"99",x"f8",x"ff",x"ff"),
   618 => (x"87",x"d6",x"02",x"a9"),
   619 => (x"89",x"c2",x"49",x"70"),
   620 => (x"bf",x"d8",x"db",x"c2"),
   621 => (x"f8",x"df",x"c2",x"91"),
   622 => (x"80",x"71",x"48",x"bf"),
   623 => (x"fc",x"58",x"a6",x"c8"),
   624 => (x"48",x"c0",x"87",x"e1"),
   625 => (x"d0",x"f0",x"8e",x"f4"),
   626 => (x"1e",x"73",x"1e",x"87"),
   627 => (x"49",x"6a",x"4a",x"71"),
   628 => (x"7a",x"71",x"81",x"c1"),
   629 => (x"bf",x"dc",x"db",x"c2"),
   630 => (x"87",x"cb",x"05",x"99"),
   631 => (x"6b",x"4b",x"a2",x"c8"),
   632 => (x"87",x"fd",x"f9",x"49"),
   633 => (x"c1",x"7b",x"49",x"70"),
   634 => (x"87",x"f1",x"ef",x"48"),
   635 => (x"71",x"1e",x"73",x"1e"),
   636 => (x"f8",x"df",x"c2",x"4b"),
   637 => (x"a3",x"c8",x"49",x"bf"),
   638 => (x"c2",x"4a",x"6a",x"4a"),
   639 => (x"d8",x"db",x"c2",x"8a"),
   640 => (x"a1",x"72",x"92",x"bf"),
   641 => (x"dc",x"db",x"c2",x"49"),
   642 => (x"9a",x"6b",x"4a",x"bf"),
   643 => (x"c8",x"49",x"a1",x"72"),
   644 => (x"e8",x"71",x"1e",x"66"),
   645 => (x"86",x"c4",x"87",x"fd"),
   646 => (x"c4",x"05",x"98",x"70"),
   647 => (x"c2",x"48",x"c0",x"87"),
   648 => (x"ee",x"48",x"c1",x"87"),
   649 => (x"5e",x"0e",x"87",x"f7"),
   650 => (x"71",x"0e",x"5c",x"5b"),
   651 => (x"72",x"4b",x"c0",x"4a"),
   652 => (x"e0",x"c0",x"02",x"9a"),
   653 => (x"49",x"a2",x"da",x"87"),
   654 => (x"c2",x"4b",x"69",x"9f"),
   655 => (x"02",x"bf",x"e0",x"db"),
   656 => (x"a2",x"d4",x"87",x"cf"),
   657 => (x"49",x"69",x"9f",x"49"),
   658 => (x"ff",x"ff",x"c0",x"4c"),
   659 => (x"c2",x"34",x"d0",x"9c"),
   660 => (x"74",x"4c",x"c0",x"87"),
   661 => (x"02",x"9b",x"73",x"b3"),
   662 => (x"c2",x"4a",x"87",x"df"),
   663 => (x"d8",x"db",x"c2",x"8a"),
   664 => (x"c2",x"92",x"49",x"bf"),
   665 => (x"48",x"bf",x"f8",x"df"),
   666 => (x"e0",x"c2",x"80",x"72"),
   667 => (x"48",x"71",x"58",x"d8"),
   668 => (x"db",x"c2",x"30",x"c4"),
   669 => (x"e9",x"c0",x"58",x"e8"),
   670 => (x"fc",x"df",x"c2",x"87"),
   671 => (x"e0",x"c2",x"4b",x"bf"),
   672 => (x"e0",x"c2",x"48",x"d4"),
   673 => (x"c2",x"78",x"bf",x"c0"),
   674 => (x"02",x"bf",x"e0",x"db"),
   675 => (x"db",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"d8"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"c4",x"e0"),
   679 => (x"db",x"c2",x"31",x"c4"),
   680 => (x"e0",x"c2",x"59",x"e8"),
   681 => (x"f2",x"ec",x"5b",x"d4"),
   682 => (x"5b",x"5e",x"0e",x"87"),
   683 => (x"f4",x"0e",x"5d",x"5c"),
   684 => (x"9a",x"4a",x"71",x"86"),
   685 => (x"c2",x"87",x"de",x"02"),
   686 => (x"c0",x"48",x"d4",x"d3"),
   687 => (x"cc",x"d3",x"c2",x"78"),
   688 => (x"d4",x"e0",x"c2",x"48"),
   689 => (x"d3",x"c2",x"78",x"bf"),
   690 => (x"e0",x"c2",x"48",x"d0"),
   691 => (x"c0",x"78",x"bf",x"d0"),
   692 => (x"c0",x"48",x"ff",x"f1"),
   693 => (x"e4",x"db",x"c2",x"78"),
   694 => (x"d3",x"c2",x"49",x"bf"),
   695 => (x"71",x"4a",x"bf",x"d4"),
   696 => (x"cb",x"c4",x"03",x"aa"),
   697 => (x"cf",x"49",x"72",x"87"),
   698 => (x"e0",x"c0",x"05",x"99"),
   699 => (x"d8",x"d3",x"c2",x"87"),
   700 => (x"cc",x"d3",x"c2",x"1e"),
   701 => (x"d3",x"c2",x"49",x"bf"),
   702 => (x"a1",x"c1",x"48",x"cc"),
   703 => (x"d2",x"e5",x"71",x"78"),
   704 => (x"c0",x"86",x"c4",x"87"),
   705 => (x"c2",x"48",x"fb",x"f1"),
   706 => (x"cc",x"78",x"d8",x"d3"),
   707 => (x"fb",x"f1",x"c0",x"87"),
   708 => (x"e0",x"c0",x"48",x"bf"),
   709 => (x"ff",x"f1",x"c0",x"80"),
   710 => (x"d4",x"d3",x"c2",x"58"),
   711 => (x"80",x"c1",x"48",x"bf"),
   712 => (x"58",x"d8",x"d3",x"c2"),
   713 => (x"00",x"0c",x"7b",x"27"),
   714 => (x"bf",x"97",x"bf",x"00"),
   715 => (x"c2",x"02",x"9c",x"4c"),
   716 => (x"e5",x"c3",x"87",x"ee"),
   717 => (x"e7",x"c2",x"02",x"ac"),
   718 => (x"fb",x"f1",x"c0",x"87"),
   719 => (x"a3",x"cb",x"4b",x"bf"),
   720 => (x"cf",x"4d",x"11",x"49"),
   721 => (x"d6",x"c1",x"05",x"ad"),
   722 => (x"df",x"49",x"74",x"87"),
   723 => (x"cd",x"89",x"c1",x"99"),
   724 => (x"e8",x"db",x"c2",x"91"),
   725 => (x"4a",x"a3",x"c1",x"81"),
   726 => (x"a3",x"c3",x"51",x"12"),
   727 => (x"c5",x"51",x"12",x"4a"),
   728 => (x"51",x"12",x"4a",x"a3"),
   729 => (x"12",x"4a",x"a3",x"c7"),
   730 => (x"4a",x"a3",x"c9",x"51"),
   731 => (x"a3",x"ce",x"51",x"12"),
   732 => (x"d0",x"51",x"12",x"4a"),
   733 => (x"51",x"12",x"4a",x"a3"),
   734 => (x"12",x"4a",x"a3",x"d2"),
   735 => (x"4a",x"a3",x"d4",x"51"),
   736 => (x"a3",x"d6",x"51",x"12"),
   737 => (x"d8",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"dc"),
   740 => (x"4a",x"a3",x"de",x"51"),
   741 => (x"f1",x"c0",x"51",x"12"),
   742 => (x"78",x"c1",x"48",x"ff"),
   743 => (x"75",x"87",x"c1",x"c1"),
   744 => (x"05",x"99",x"c8",x"49"),
   745 => (x"75",x"87",x"f3",x"c0"),
   746 => (x"05",x"99",x"d0",x"49"),
   747 => (x"66",x"dc",x"87",x"d0"),
   748 => (x"87",x"ca",x"c0",x"02"),
   749 => (x"66",x"dc",x"49",x"73"),
   750 => (x"02",x"98",x"70",x"0f"),
   751 => (x"f1",x"c0",x"87",x"dc"),
   752 => (x"c0",x"05",x"bf",x"ff"),
   753 => (x"db",x"c2",x"87",x"c6"),
   754 => (x"50",x"c0",x"48",x"e8"),
   755 => (x"48",x"ff",x"f1",x"c0"),
   756 => (x"f1",x"c0",x"78",x"c0"),
   757 => (x"c2",x"48",x"bf",x"fb"),
   758 => (x"f1",x"c0",x"87",x"dc"),
   759 => (x"78",x"c0",x"48",x"ff"),
   760 => (x"bf",x"e4",x"db",x"c2"),
   761 => (x"d4",x"d3",x"c2",x"49"),
   762 => (x"aa",x"71",x"4a",x"bf"),
   763 => (x"87",x"f5",x"fb",x"04"),
   764 => (x"bf",x"d4",x"e0",x"c2"),
   765 => (x"87",x"c8",x"c0",x"05"),
   766 => (x"bf",x"e0",x"db",x"c2"),
   767 => (x"87",x"f4",x"c1",x"02"),
   768 => (x"bf",x"d0",x"d3",x"c2"),
   769 => (x"87",x"d9",x"f1",x"49"),
   770 => (x"58",x"d4",x"d3",x"c2"),
   771 => (x"db",x"c2",x"7e",x"70"),
   772 => (x"c0",x"02",x"bf",x"e0"),
   773 => (x"49",x"6e",x"87",x"dd"),
   774 => (x"ff",x"ff",x"ff",x"cf"),
   775 => (x"02",x"a9",x"99",x"f8"),
   776 => (x"c4",x"87",x"c8",x"c0"),
   777 => (x"78",x"c0",x"48",x"a6"),
   778 => (x"c4",x"87",x"e6",x"c0"),
   779 => (x"78",x"c1",x"48",x"a6"),
   780 => (x"6e",x"87",x"de",x"c0"),
   781 => (x"f8",x"ff",x"cf",x"49"),
   782 => (x"c0",x"02",x"a9",x"99"),
   783 => (x"a6",x"c8",x"87",x"c8"),
   784 => (x"c0",x"78",x"c0",x"48"),
   785 => (x"a6",x"c8",x"87",x"c5"),
   786 => (x"c4",x"78",x"c1",x"48"),
   787 => (x"66",x"c8",x"48",x"a6"),
   788 => (x"05",x"66",x"c4",x"78"),
   789 => (x"6e",x"87",x"dd",x"c0"),
   790 => (x"c2",x"89",x"c2",x"49"),
   791 => (x"91",x"bf",x"d8",x"db"),
   792 => (x"bf",x"f8",x"df",x"c2"),
   793 => (x"c2",x"80",x"71",x"48"),
   794 => (x"c2",x"58",x"d0",x"d3"),
   795 => (x"c0",x"48",x"d4",x"d3"),
   796 => (x"87",x"e1",x"f9",x"78"),
   797 => (x"8e",x"f4",x"48",x"c0"),
   798 => (x"00",x"87",x"de",x"e5"),
   799 => (x"00",x"00",x"00",x"00"),
   800 => (x"1e",x"00",x"00",x"00"),
   801 => (x"c3",x"48",x"d4",x"ff"),
   802 => (x"49",x"68",x"78",x"ff"),
   803 => (x"87",x"c6",x"02",x"99"),
   804 => (x"05",x"a9",x"fb",x"c0"),
   805 => (x"48",x"71",x"87",x"ee"),
   806 => (x"5e",x"0e",x"4f",x"26"),
   807 => (x"71",x"0e",x"5c",x"5b"),
   808 => (x"ff",x"4b",x"c0",x"4a"),
   809 => (x"ff",x"c3",x"48",x"d4"),
   810 => (x"99",x"49",x"68",x"78"),
   811 => (x"87",x"c1",x"c1",x"02"),
   812 => (x"02",x"a9",x"ec",x"c0"),
   813 => (x"c0",x"87",x"fa",x"c0"),
   814 => (x"c0",x"02",x"a9",x"fb"),
   815 => (x"66",x"cc",x"87",x"f3"),
   816 => (x"cc",x"03",x"ab",x"b7"),
   817 => (x"02",x"66",x"d0",x"87"),
   818 => (x"09",x"72",x"87",x"c7"),
   819 => (x"c1",x"09",x"79",x"97"),
   820 => (x"02",x"99",x"71",x"82"),
   821 => (x"83",x"c1",x"87",x"c2"),
   822 => (x"c3",x"48",x"d4",x"ff"),
   823 => (x"49",x"68",x"78",x"ff"),
   824 => (x"87",x"cd",x"02",x"99"),
   825 => (x"02",x"a9",x"ec",x"c0"),
   826 => (x"fb",x"c0",x"87",x"c7"),
   827 => (x"cd",x"ff",x"05",x"a9"),
   828 => (x"02",x"66",x"d0",x"87"),
   829 => (x"97",x"c0",x"87",x"c3"),
   830 => (x"a9",x"fb",x"c0",x"7a"),
   831 => (x"73",x"87",x"c7",x"05"),
   832 => (x"8c",x"0c",x"c0",x"4c"),
   833 => (x"4c",x"73",x"87",x"c2"),
   834 => (x"87",x"c2",x"48",x"74"),
   835 => (x"4c",x"26",x"4d",x"26"),
   836 => (x"4f",x"26",x"4b",x"26"),
   837 => (x"48",x"d4",x"ff",x"1e"),
   838 => (x"68",x"78",x"ff",x"c3"),
   839 => (x"b7",x"f0",x"c0",x"49"),
   840 => (x"87",x"ca",x"04",x"a9"),
   841 => (x"a9",x"b7",x"f9",x"c0"),
   842 => (x"c0",x"87",x"c3",x"01"),
   843 => (x"c1",x"c1",x"89",x"f0"),
   844 => (x"ca",x"04",x"a9",x"b7"),
   845 => (x"b7",x"c6",x"c1",x"87"),
   846 => (x"87",x"c3",x"01",x"a9"),
   847 => (x"71",x"89",x"f7",x"c0"),
   848 => (x"0e",x"4f",x"26",x"48"),
   849 => (x"5d",x"5c",x"5b",x"5e"),
   850 => (x"71",x"86",x"f4",x"0e"),
   851 => (x"4b",x"d4",x"ff",x"4c"),
   852 => (x"c3",x"7e",x"4d",x"c0"),
   853 => (x"d0",x"ff",x"7b",x"ff"),
   854 => (x"c0",x"c8",x"48",x"bf"),
   855 => (x"a6",x"c8",x"98",x"c0"),
   856 => (x"02",x"98",x"70",x"58"),
   857 => (x"d0",x"ff",x"87",x"d0"),
   858 => (x"c0",x"c8",x"48",x"bf"),
   859 => (x"a6",x"c8",x"98",x"c0"),
   860 => (x"05",x"98",x"70",x"58"),
   861 => (x"d0",x"ff",x"87",x"f0"),
   862 => (x"78",x"e1",x"c0",x"48"),
   863 => (x"c2",x"fc",x"7b",x"d4"),
   864 => (x"99",x"49",x"70",x"87"),
   865 => (x"87",x"c7",x"c1",x"02"),
   866 => (x"c8",x"7b",x"ff",x"c3"),
   867 => (x"78",x"6b",x"48",x"a6"),
   868 => (x"c0",x"48",x"66",x"c8"),
   869 => (x"c8",x"02",x"a8",x"fb"),
   870 => (x"f0",x"e0",x"c2",x"87"),
   871 => (x"ee",x"c0",x"02",x"bf"),
   872 => (x"71",x"4d",x"c1",x"87"),
   873 => (x"e6",x"c0",x"02",x"99"),
   874 => (x"a9",x"fb",x"c0",x"87"),
   875 => (x"fb",x"87",x"c3",x"02"),
   876 => (x"ff",x"c3",x"87",x"d1"),
   877 => (x"c1",x"49",x"6b",x"7b"),
   878 => (x"cc",x"05",x"a9",x"c6"),
   879 => (x"7b",x"ff",x"c3",x"87"),
   880 => (x"48",x"a6",x"c8",x"7b"),
   881 => (x"49",x"c0",x"78",x"6b"),
   882 => (x"05",x"99",x"71",x"4d"),
   883 => (x"75",x"87",x"da",x"ff"),
   884 => (x"de",x"c1",x"05",x"9d"),
   885 => (x"7b",x"ff",x"c3",x"87"),
   886 => (x"ff",x"c3",x"4a",x"6b"),
   887 => (x"48",x"a6",x"c4",x"7b"),
   888 => (x"48",x"6e",x"78",x"6b"),
   889 => (x"a6",x"c4",x"80",x"c1"),
   890 => (x"49",x"a4",x"c8",x"58"),
   891 => (x"c8",x"49",x"69",x"97"),
   892 => (x"da",x"05",x"a9",x"66"),
   893 => (x"49",x"a4",x"c9",x"87"),
   894 => (x"aa",x"49",x"69",x"97"),
   895 => (x"ca",x"87",x"d0",x"05"),
   896 => (x"69",x"97",x"49",x"a4"),
   897 => (x"a9",x"66",x"c4",x"49"),
   898 => (x"c1",x"87",x"c4",x"05"),
   899 => (x"c8",x"87",x"d6",x"4d"),
   900 => (x"ec",x"c0",x"48",x"66"),
   901 => (x"87",x"c9",x"02",x"a8"),
   902 => (x"c0",x"48",x"66",x"c8"),
   903 => (x"c4",x"05",x"a8",x"fb"),
   904 => (x"c1",x"7e",x"c0",x"87"),
   905 => (x"7b",x"ff",x"c3",x"4d"),
   906 => (x"6b",x"48",x"a6",x"c8"),
   907 => (x"02",x"9d",x"75",x"78"),
   908 => (x"ff",x"87",x"e2",x"fe"),
   909 => (x"c8",x"48",x"bf",x"d0"),
   910 => (x"c8",x"98",x"c0",x"c0"),
   911 => (x"98",x"70",x"58",x"a6"),
   912 => (x"ff",x"87",x"d0",x"02"),
   913 => (x"c8",x"48",x"bf",x"d0"),
   914 => (x"c8",x"98",x"c0",x"c0"),
   915 => (x"98",x"70",x"58",x"a6"),
   916 => (x"ff",x"87",x"f0",x"05"),
   917 => (x"e0",x"c0",x"48",x"d0"),
   918 => (x"f4",x"48",x"6e",x"78"),
   919 => (x"87",x"ec",x"fa",x"8e"),
   920 => (x"5c",x"5b",x"5e",x"0e"),
   921 => (x"86",x"f4",x"0e",x"5d"),
   922 => (x"ff",x"59",x"a6",x"c4"),
   923 => (x"c0",x"c8",x"4c",x"d0"),
   924 => (x"1e",x"6e",x"4b",x"c0"),
   925 => (x"49",x"f4",x"e0",x"c2"),
   926 => (x"c4",x"87",x"cf",x"e9"),
   927 => (x"02",x"98",x"70",x"86"),
   928 => (x"c2",x"87",x"f7",x"c5"),
   929 => (x"4d",x"bf",x"f8",x"e0"),
   930 => (x"f6",x"fa",x"49",x"6e"),
   931 => (x"58",x"a6",x"c8",x"87"),
   932 => (x"98",x"73",x"48",x"6c"),
   933 => (x"70",x"58",x"a6",x"cc"),
   934 => (x"87",x"cc",x"02",x"98"),
   935 => (x"98",x"73",x"48",x"6c"),
   936 => (x"70",x"58",x"a6",x"c4"),
   937 => (x"87",x"f4",x"05",x"98"),
   938 => (x"d4",x"ff",x"7c",x"c5"),
   939 => (x"78",x"d5",x"c1",x"48"),
   940 => (x"bf",x"f0",x"e0",x"c2"),
   941 => (x"c4",x"81",x"c1",x"49"),
   942 => (x"8a",x"c1",x"4a",x"66"),
   943 => (x"48",x"72",x"32",x"c6"),
   944 => (x"d4",x"ff",x"b0",x"71"),
   945 => (x"48",x"6c",x"78",x"08"),
   946 => (x"a6",x"c4",x"98",x"73"),
   947 => (x"02",x"98",x"70",x"58"),
   948 => (x"48",x"6c",x"87",x"cc"),
   949 => (x"a6",x"c4",x"98",x"73"),
   950 => (x"05",x"98",x"70",x"58"),
   951 => (x"7c",x"c4",x"87",x"f4"),
   952 => (x"c3",x"48",x"d4",x"ff"),
   953 => (x"48",x"6c",x"78",x"ff"),
   954 => (x"a6",x"c4",x"98",x"73"),
   955 => (x"02",x"98",x"70",x"58"),
   956 => (x"48",x"6c",x"87",x"cc"),
   957 => (x"a6",x"c4",x"98",x"73"),
   958 => (x"05",x"98",x"70",x"58"),
   959 => (x"7c",x"c5",x"87",x"f4"),
   960 => (x"c1",x"48",x"d4",x"ff"),
   961 => (x"78",x"c1",x"78",x"d3"),
   962 => (x"98",x"73",x"48",x"6c"),
   963 => (x"70",x"58",x"a6",x"c4"),
   964 => (x"87",x"cc",x"02",x"98"),
   965 => (x"98",x"73",x"48",x"6c"),
   966 => (x"70",x"58",x"a6",x"c4"),
   967 => (x"87",x"f4",x"05",x"98"),
   968 => (x"9d",x"75",x"7c",x"c4"),
   969 => (x"87",x"d0",x"c2",x"02"),
   970 => (x"7e",x"d8",x"d3",x"c2"),
   971 => (x"f4",x"e0",x"c2",x"1e"),
   972 => (x"87",x"f8",x"ea",x"49"),
   973 => (x"98",x"70",x"86",x"c4"),
   974 => (x"c0",x"87",x"c5",x"05"),
   975 => (x"87",x"fc",x"c2",x"48"),
   976 => (x"ad",x"b7",x"c0",x"c8"),
   977 => (x"4a",x"87",x"c4",x"04"),
   978 => (x"75",x"87",x"c4",x"8d"),
   979 => (x"6c",x"4d",x"c0",x"4a"),
   980 => (x"c8",x"98",x"73",x"48"),
   981 => (x"98",x"70",x"58",x"a6"),
   982 => (x"6c",x"87",x"cc",x"02"),
   983 => (x"c8",x"98",x"73",x"48"),
   984 => (x"98",x"70",x"58",x"a6"),
   985 => (x"cd",x"87",x"f4",x"05"),
   986 => (x"48",x"d4",x"ff",x"7c"),
   987 => (x"72",x"78",x"d4",x"c1"),
   988 => (x"71",x"8a",x"c1",x"49"),
   989 => (x"87",x"d9",x"02",x"99"),
   990 => (x"48",x"bf",x"97",x"6e"),
   991 => (x"78",x"08",x"d4",x"ff"),
   992 => (x"80",x"c1",x"48",x"6e"),
   993 => (x"72",x"58",x"a6",x"c4"),
   994 => (x"71",x"8a",x"c1",x"49"),
   995 => (x"e7",x"ff",x"05",x"99"),
   996 => (x"73",x"48",x"6c",x"87"),
   997 => (x"58",x"a6",x"c4",x"98"),
   998 => (x"cc",x"02",x"98",x"70"),
   999 => (x"73",x"48",x"6c",x"87"),
  1000 => (x"58",x"a6",x"c4",x"98"),
  1001 => (x"f4",x"05",x"98",x"70"),
  1002 => (x"c2",x"7c",x"c4",x"87"),
  1003 => (x"e8",x"49",x"f4",x"e0"),
  1004 => (x"9d",x"75",x"87",x"d7"),
  1005 => (x"87",x"f0",x"fd",x"05"),
  1006 => (x"98",x"73",x"48",x"6c"),
  1007 => (x"70",x"58",x"a6",x"c4"),
  1008 => (x"87",x"cd",x"02",x"98"),
  1009 => (x"98",x"73",x"48",x"6c"),
  1010 => (x"70",x"58",x"a6",x"c4"),
  1011 => (x"f3",x"ff",x"05",x"98"),
  1012 => (x"ff",x"7c",x"c5",x"87"),
  1013 => (x"d3",x"c1",x"48",x"d4"),
  1014 => (x"6c",x"78",x"c0",x"78"),
  1015 => (x"c4",x"98",x"73",x"48"),
  1016 => (x"98",x"70",x"58",x"a6"),
  1017 => (x"6c",x"87",x"cd",x"02"),
  1018 => (x"c4",x"98",x"73",x"48"),
  1019 => (x"98",x"70",x"58",x"a6"),
  1020 => (x"87",x"f3",x"ff",x"05"),
  1021 => (x"48",x"c1",x"7c",x"c4"),
  1022 => (x"48",x"c0",x"87",x"c2"),
  1023 => (x"cb",x"f4",x"8e",x"f4"),
  1024 => (x"5b",x"5e",x"0e",x"87"),
  1025 => (x"1e",x"0e",x"5d",x"5c"),
  1026 => (x"4c",x"c0",x"4b",x"71"),
  1027 => (x"04",x"ab",x"b7",x"4d"),
  1028 => (x"c0",x"87",x"e9",x"c0"),
  1029 => (x"75",x"1e",x"c3",x"f5"),
  1030 => (x"87",x"c4",x"02",x"9d"),
  1031 => (x"87",x"c2",x"4a",x"c0"),
  1032 => (x"49",x"72",x"4a",x"c1"),
  1033 => (x"c4",x"87",x"c2",x"ea"),
  1034 => (x"c1",x"58",x"a6",x"86"),
  1035 => (x"c2",x"05",x"6e",x"84"),
  1036 => (x"c1",x"4c",x"73",x"87"),
  1037 => (x"ac",x"b7",x"73",x"85"),
  1038 => (x"87",x"d7",x"ff",x"06"),
  1039 => (x"f3",x"26",x"48",x"6e"),
  1040 => (x"5e",x"0e",x"87",x"ca"),
  1041 => (x"0e",x"5d",x"5c",x"5b"),
  1042 => (x"49",x"4c",x"71",x"1e"),
  1043 => (x"bf",x"c4",x"e1",x"c2"),
  1044 => (x"87",x"ed",x"fe",x"81"),
  1045 => (x"02",x"9d",x"4d",x"70"),
  1046 => (x"c2",x"87",x"fc",x"c0"),
  1047 => (x"75",x"4b",x"e8",x"db"),
  1048 => (x"ff",x"49",x"cb",x"4a"),
  1049 => (x"74",x"87",x"c9",x"c1"),
  1050 => (x"c2",x"91",x"de",x"49"),
  1051 => (x"71",x"48",x"d8",x"e1"),
  1052 => (x"58",x"a6",x"c4",x"80"),
  1053 => (x"48",x"e7",x"c2",x"c1"),
  1054 => (x"a1",x"c8",x"49",x"6e"),
  1055 => (x"71",x"41",x"20",x"4a"),
  1056 => (x"87",x"f9",x"05",x"aa"),
  1057 => (x"51",x"10",x"51",x"10"),
  1058 => (x"49",x"74",x"51",x"10"),
  1059 => (x"87",x"fd",x"c4",x"c1"),
  1060 => (x"49",x"e8",x"db",x"c2"),
  1061 => (x"c1",x"87",x"c9",x"f7"),
  1062 => (x"c1",x"49",x"f8",x"e3"),
  1063 => (x"c1",x"87",x"c0",x"c6"),
  1064 => (x"26",x"87",x"cf",x"c6"),
  1065 => (x"4c",x"87",x"e5",x"f1"),
  1066 => (x"69",x"64",x"61",x"6f"),
  1067 => (x"2e",x"2e",x"67",x"6e"),
  1068 => (x"20",x"80",x"00",x"2e"),
  1069 => (x"6b",x"63",x"61",x"42"),
  1070 => (x"61",x"6f",x"4c",x"00"),
  1071 => (x"2e",x"2a",x"20",x"64"),
  1072 => (x"20",x"3a",x"00",x"20"),
  1073 => (x"42",x"20",x"80",x"00"),
  1074 => (x"00",x"6b",x"63",x"61"),
  1075 => (x"78",x"45",x"20",x"80"),
  1076 => (x"53",x"00",x"74",x"69"),
  1077 => (x"6e",x"49",x"20",x"44"),
  1078 => (x"2e",x"2e",x"74",x"69"),
  1079 => (x"00",x"4b",x"4f",x"00"),
  1080 => (x"54",x"4f",x"4f",x"42"),
  1081 => (x"20",x"20",x"20",x"20"),
  1082 => (x"00",x"4d",x"4f",x"52"),
  1083 => (x"71",x"1e",x"73",x"1e"),
  1084 => (x"e1",x"c2",x"49",x"4b"),
  1085 => (x"fc",x"81",x"bf",x"c4"),
  1086 => (x"4a",x"70",x"87",x"c7"),
  1087 => (x"87",x"c4",x"02",x"9a"),
  1088 => (x"87",x"e2",x"e4",x"49"),
  1089 => (x"48",x"c4",x"e1",x"c2"),
  1090 => (x"49",x"73",x"78",x"c0"),
  1091 => (x"ef",x"87",x"e9",x"c1"),
  1092 => (x"73",x"1e",x"87",x"fe"),
  1093 => (x"c4",x"4b",x"71",x"1e"),
  1094 => (x"c1",x"02",x"4a",x"a3"),
  1095 => (x"8a",x"c1",x"87",x"c8"),
  1096 => (x"8a",x"87",x"dc",x"02"),
  1097 => (x"87",x"f1",x"c0",x"02"),
  1098 => (x"c4",x"c1",x"05",x"8a"),
  1099 => (x"c4",x"e1",x"c2",x"87"),
  1100 => (x"fc",x"c0",x"02",x"bf"),
  1101 => (x"88",x"c1",x"48",x"87"),
  1102 => (x"58",x"c8",x"e1",x"c2"),
  1103 => (x"c2",x"87",x"f2",x"c0"),
  1104 => (x"49",x"bf",x"c4",x"e1"),
  1105 => (x"e1",x"c2",x"89",x"d0"),
  1106 => (x"b7",x"c0",x"59",x"c8"),
  1107 => (x"e0",x"c0",x"03",x"a9"),
  1108 => (x"c4",x"e1",x"c2",x"87"),
  1109 => (x"d8",x"78",x"c0",x"48"),
  1110 => (x"c4",x"e1",x"c2",x"87"),
  1111 => (x"80",x"c1",x"48",x"bf"),
  1112 => (x"58",x"c8",x"e1",x"c2"),
  1113 => (x"e1",x"c2",x"87",x"cb"),
  1114 => (x"d0",x"48",x"bf",x"c4"),
  1115 => (x"c8",x"e1",x"c2",x"80"),
  1116 => (x"c3",x"49",x"73",x"58"),
  1117 => (x"87",x"d8",x"ee",x"87"),
  1118 => (x"5c",x"5b",x"5e",x"0e"),
  1119 => (x"86",x"f0",x"0e",x"5d"),
  1120 => (x"c2",x"59",x"a6",x"d0"),
  1121 => (x"c0",x"4d",x"d8",x"d3"),
  1122 => (x"48",x"a6",x"c4",x"4c"),
  1123 => (x"e1",x"c2",x"78",x"c0"),
  1124 => (x"c0",x"48",x"bf",x"c4"),
  1125 => (x"c1",x"06",x"a8",x"b7"),
  1126 => (x"d3",x"c2",x"87",x"c1"),
  1127 => (x"02",x"98",x"48",x"d8"),
  1128 => (x"c0",x"87",x"f8",x"c0"),
  1129 => (x"c8",x"1e",x"c3",x"f5"),
  1130 => (x"87",x"c7",x"02",x"66"),
  1131 => (x"c0",x"48",x"a6",x"c4"),
  1132 => (x"c4",x"87",x"c5",x"78"),
  1133 => (x"78",x"c1",x"48",x"a6"),
  1134 => (x"e3",x"49",x"66",x"c4"),
  1135 => (x"86",x"c4",x"87",x"eb"),
  1136 => (x"84",x"c1",x"4d",x"70"),
  1137 => (x"c1",x"48",x"66",x"c4"),
  1138 => (x"58",x"a6",x"c8",x"80"),
  1139 => (x"bf",x"c4",x"e1",x"c2"),
  1140 => (x"c6",x"03",x"ac",x"b7"),
  1141 => (x"05",x"9d",x"75",x"87"),
  1142 => (x"c0",x"87",x"c8",x"ff"),
  1143 => (x"02",x"9d",x"75",x"4c"),
  1144 => (x"c0",x"87",x"de",x"c3"),
  1145 => (x"c8",x"1e",x"c3",x"f5"),
  1146 => (x"87",x"c7",x"02",x"66"),
  1147 => (x"c0",x"48",x"a6",x"cc"),
  1148 => (x"cc",x"87",x"c5",x"78"),
  1149 => (x"78",x"c1",x"48",x"a6"),
  1150 => (x"e2",x"49",x"66",x"cc"),
  1151 => (x"86",x"c4",x"87",x"eb"),
  1152 => (x"02",x"6e",x"58",x"a6"),
  1153 => (x"49",x"87",x"e6",x"c2"),
  1154 => (x"69",x"97",x"81",x"cb"),
  1155 => (x"02",x"99",x"d0",x"49"),
  1156 => (x"c1",x"87",x"d6",x"c1"),
  1157 => (x"74",x"4a",x"ec",x"c3"),
  1158 => (x"c1",x"91",x"cb",x"49"),
  1159 => (x"72",x"81",x"f8",x"e3"),
  1160 => (x"c3",x"81",x"c8",x"79"),
  1161 => (x"49",x"74",x"51",x"ff"),
  1162 => (x"e1",x"c2",x"91",x"de"),
  1163 => (x"85",x"71",x"4d",x"d8"),
  1164 => (x"7d",x"97",x"c1",x"c2"),
  1165 => (x"c0",x"49",x"a5",x"c1"),
  1166 => (x"db",x"c2",x"51",x"e0"),
  1167 => (x"02",x"bf",x"97",x"e8"),
  1168 => (x"84",x"c1",x"87",x"d2"),
  1169 => (x"c2",x"4b",x"a5",x"c2"),
  1170 => (x"db",x"4a",x"e8",x"db"),
  1171 => (x"df",x"f9",x"fe",x"49"),
  1172 => (x"87",x"d9",x"c1",x"87"),
  1173 => (x"c0",x"49",x"a5",x"cd"),
  1174 => (x"c2",x"84",x"c1",x"51"),
  1175 => (x"4a",x"6e",x"4b",x"a5"),
  1176 => (x"f9",x"fe",x"49",x"cb"),
  1177 => (x"c4",x"c1",x"87",x"ca"),
  1178 => (x"cb",x"49",x"74",x"87"),
  1179 => (x"f8",x"e3",x"c1",x"91"),
  1180 => (x"c2",x"c1",x"c1",x"81"),
  1181 => (x"e8",x"db",x"c2",x"79"),
  1182 => (x"d8",x"02",x"bf",x"97"),
  1183 => (x"de",x"49",x"74",x"87"),
  1184 => (x"c2",x"84",x"c1",x"91"),
  1185 => (x"71",x"4b",x"d8",x"e1"),
  1186 => (x"e8",x"db",x"c2",x"83"),
  1187 => (x"fe",x"49",x"dd",x"4a"),
  1188 => (x"d8",x"87",x"dd",x"f8"),
  1189 => (x"de",x"4b",x"74",x"87"),
  1190 => (x"d8",x"e1",x"c2",x"93"),
  1191 => (x"49",x"a3",x"cb",x"83"),
  1192 => (x"84",x"c1",x"51",x"c0"),
  1193 => (x"cb",x"4a",x"6e",x"73"),
  1194 => (x"c3",x"f8",x"fe",x"49"),
  1195 => (x"48",x"66",x"c4",x"87"),
  1196 => (x"a6",x"c8",x"80",x"c1"),
  1197 => (x"ac",x"b7",x"c7",x"58"),
  1198 => (x"87",x"c5",x"c0",x"03"),
  1199 => (x"e2",x"fc",x"05",x"6e"),
  1200 => (x"ac",x"b7",x"c7",x"87"),
  1201 => (x"87",x"d3",x"c0",x"03"),
  1202 => (x"91",x"de",x"49",x"74"),
  1203 => (x"81",x"d8",x"e1",x"c2"),
  1204 => (x"84",x"c1",x"51",x"c0"),
  1205 => (x"04",x"ac",x"b7",x"c7"),
  1206 => (x"c1",x"87",x"ed",x"ff"),
  1207 => (x"c0",x"48",x"cd",x"e5"),
  1208 => (x"c5",x"e5",x"c1",x"50"),
  1209 => (x"d3",x"cc",x"c1",x"48"),
  1210 => (x"c9",x"e5",x"c1",x"78"),
  1211 => (x"f2",x"c2",x"c1",x"48"),
  1212 => (x"d0",x"e5",x"c1",x"78"),
  1213 => (x"d2",x"c4",x"c1",x"48"),
  1214 => (x"49",x"66",x"cc",x"78"),
  1215 => (x"87",x"cd",x"fb",x"c0"),
  1216 => (x"c7",x"e8",x"8e",x"f0"),
  1217 => (x"4a",x"71",x"1e",x"87"),
  1218 => (x"5a",x"f4",x"e0",x"c2"),
  1219 => (x"e7",x"f9",x"49",x"72"),
  1220 => (x"1e",x"4f",x"26",x"87"),
  1221 => (x"cb",x"49",x"4a",x"71"),
  1222 => (x"f8",x"e3",x"c1",x"91"),
  1223 => (x"11",x"81",x"c8",x"81"),
  1224 => (x"f0",x"e0",x"c2",x"48"),
  1225 => (x"a2",x"f0",x"c0",x"58"),
  1226 => (x"d3",x"f6",x"fe",x"49"),
  1227 => (x"d5",x"49",x"c0",x"87"),
  1228 => (x"4f",x"26",x"87",x"c0"),
  1229 => (x"5c",x"5b",x"5e",x"0e"),
  1230 => (x"86",x"f0",x"0e",x"5d"),
  1231 => (x"cb",x"49",x"4d",x"71"),
  1232 => (x"f8",x"e3",x"c1",x"91"),
  1233 => (x"7e",x"a1",x"ca",x"81"),
  1234 => (x"c2",x"48",x"a6",x"c4"),
  1235 => (x"78",x"bf",x"e8",x"e0"),
  1236 => (x"4a",x"bf",x"97",x"6e"),
  1237 => (x"72",x"4b",x"66",x"c4"),
  1238 => (x"4a",x"a1",x"c8",x"2b"),
  1239 => (x"a6",x"cc",x"48",x"12"),
  1240 => (x"c1",x"9b",x"70",x"58"),
  1241 => (x"97",x"81",x"c9",x"83"),
  1242 => (x"ab",x"b7",x"49",x"69"),
  1243 => (x"c0",x"87",x"c2",x"04"),
  1244 => (x"bf",x"97",x"6e",x"4b"),
  1245 => (x"49",x"66",x"c8",x"4a"),
  1246 => (x"b9",x"ff",x"31",x"72"),
  1247 => (x"73",x"99",x"66",x"c4"),
  1248 => (x"71",x"34",x"72",x"4c"),
  1249 => (x"ec",x"e0",x"c2",x"b4"),
  1250 => (x"48",x"d4",x"ff",x"5c"),
  1251 => (x"ff",x"78",x"ff",x"c3"),
  1252 => (x"c8",x"48",x"bf",x"d0"),
  1253 => (x"d0",x"98",x"c0",x"c0"),
  1254 => (x"98",x"70",x"58",x"a6"),
  1255 => (x"ff",x"87",x"d0",x"02"),
  1256 => (x"c8",x"48",x"bf",x"d0"),
  1257 => (x"c4",x"98",x"c0",x"c0"),
  1258 => (x"98",x"70",x"58",x"a6"),
  1259 => (x"ff",x"87",x"f0",x"05"),
  1260 => (x"e1",x"c0",x"48",x"d0"),
  1261 => (x"48",x"d4",x"ff",x"78"),
  1262 => (x"0c",x"70",x"78",x"de"),
  1263 => (x"48",x"74",x"0c",x"7c"),
  1264 => (x"ff",x"28",x"b7",x"c8"),
  1265 => (x"74",x"78",x"08",x"d4"),
  1266 => (x"28",x"b7",x"d0",x"48"),
  1267 => (x"78",x"08",x"d4",x"ff"),
  1268 => (x"b7",x"d8",x"48",x"74"),
  1269 => (x"08",x"d4",x"ff",x"28"),
  1270 => (x"bf",x"d0",x"ff",x"78"),
  1271 => (x"c0",x"c0",x"c8",x"48"),
  1272 => (x"58",x"a6",x"c4",x"98"),
  1273 => (x"d0",x"02",x"98",x"70"),
  1274 => (x"bf",x"d0",x"ff",x"87"),
  1275 => (x"c0",x"c0",x"c8",x"48"),
  1276 => (x"58",x"a6",x"c4",x"98"),
  1277 => (x"f0",x"05",x"98",x"70"),
  1278 => (x"48",x"d0",x"ff",x"87"),
  1279 => (x"c7",x"78",x"e0",x"c0"),
  1280 => (x"c1",x"1e",x"c0",x"1e"),
  1281 => (x"c2",x"1e",x"f8",x"e3"),
  1282 => (x"49",x"bf",x"ec",x"e0"),
  1283 => (x"75",x"87",x"e1",x"c1"),
  1284 => (x"f8",x"f6",x"c0",x"49"),
  1285 => (x"e3",x"8e",x"e4",x"87"),
  1286 => (x"73",x"1e",x"87",x"f2"),
  1287 => (x"49",x"4b",x"71",x"1e"),
  1288 => (x"73",x"87",x"d1",x"fc"),
  1289 => (x"87",x"cc",x"fc",x"49"),
  1290 => (x"1e",x"87",x"e5",x"e3"),
  1291 => (x"4b",x"71",x"1e",x"73"),
  1292 => (x"02",x"4a",x"a3",x"c2"),
  1293 => (x"8a",x"c1",x"87",x"d5"),
  1294 => (x"c2",x"87",x"db",x"05"),
  1295 => (x"02",x"bf",x"c0",x"e1"),
  1296 => (x"c1",x"48",x"87",x"d4"),
  1297 => (x"c4",x"e1",x"c2",x"88"),
  1298 => (x"c2",x"87",x"cb",x"58"),
  1299 => (x"48",x"bf",x"c0",x"e1"),
  1300 => (x"e1",x"c2",x"80",x"c1"),
  1301 => (x"1e",x"c7",x"58",x"c4"),
  1302 => (x"e3",x"c1",x"1e",x"c0"),
  1303 => (x"e0",x"c2",x"1e",x"f8"),
  1304 => (x"cb",x"49",x"bf",x"ec"),
  1305 => (x"c0",x"49",x"73",x"87"),
  1306 => (x"f4",x"87",x"e2",x"f5"),
  1307 => (x"87",x"e0",x"e2",x"8e"),
  1308 => (x"5c",x"5b",x"5e",x"0e"),
  1309 => (x"d8",x"ff",x"0e",x"5d"),
  1310 => (x"59",x"a6",x"dc",x"86"),
  1311 => (x"c0",x"48",x"a6",x"c8"),
  1312 => (x"c0",x"80",x"c4",x"78"),
  1313 => (x"80",x"c4",x"4d",x"78"),
  1314 => (x"bf",x"c0",x"e1",x"c2"),
  1315 => (x"48",x"d4",x"ff",x"78"),
  1316 => (x"ff",x"78",x"ff",x"c3"),
  1317 => (x"c8",x"48",x"bf",x"d0"),
  1318 => (x"c4",x"98",x"c0",x"c0"),
  1319 => (x"98",x"70",x"58",x"a6"),
  1320 => (x"ff",x"87",x"d0",x"02"),
  1321 => (x"c8",x"48",x"bf",x"d0"),
  1322 => (x"c4",x"98",x"c0",x"c0"),
  1323 => (x"98",x"70",x"58",x"a6"),
  1324 => (x"ff",x"87",x"f0",x"05"),
  1325 => (x"e1",x"c0",x"48",x"d0"),
  1326 => (x"48",x"d4",x"ff",x"78"),
  1327 => (x"df",x"ff",x"78",x"d4"),
  1328 => (x"d4",x"ff",x"87",x"c1"),
  1329 => (x"78",x"ff",x"c3",x"48"),
  1330 => (x"ff",x"48",x"a6",x"d4"),
  1331 => (x"d4",x"78",x"bf",x"d4"),
  1332 => (x"fb",x"c0",x"48",x"66"),
  1333 => (x"d1",x"c1",x"02",x"a8"),
  1334 => (x"66",x"f8",x"c0",x"87"),
  1335 => (x"6a",x"82",x"c4",x"4a"),
  1336 => (x"c1",x"1e",x"72",x"7e"),
  1337 => (x"c4",x"48",x"f9",x"c2"),
  1338 => (x"a1",x"c8",x"49",x"66"),
  1339 => (x"71",x"41",x"20",x"4a"),
  1340 => (x"87",x"f9",x"05",x"aa"),
  1341 => (x"4a",x"26",x"51",x"10"),
  1342 => (x"48",x"66",x"f8",x"c0"),
  1343 => (x"78",x"c5",x"cc",x"c1"),
  1344 => (x"81",x"c7",x"49",x"6a"),
  1345 => (x"c1",x"51",x"66",x"d4"),
  1346 => (x"6a",x"1e",x"d8",x"1e"),
  1347 => (x"ff",x"81",x"c8",x"49"),
  1348 => (x"c8",x"87",x"c7",x"de"),
  1349 => (x"48",x"66",x"d0",x"86"),
  1350 => (x"01",x"a8",x"b7",x"c0"),
  1351 => (x"4d",x"c1",x"87",x"c4"),
  1352 => (x"66",x"d0",x"87",x"c8"),
  1353 => (x"d4",x"88",x"c1",x"48"),
  1354 => (x"66",x"d4",x"58",x"a6"),
  1355 => (x"87",x"e5",x"ca",x"02"),
  1356 => (x"b7",x"66",x"c0",x"c1"),
  1357 => (x"dc",x"ca",x"03",x"ad"),
  1358 => (x"48",x"d4",x"ff",x"87"),
  1359 => (x"d4",x"78",x"ff",x"c3"),
  1360 => (x"d4",x"ff",x"48",x"a6"),
  1361 => (x"66",x"d4",x"78",x"bf"),
  1362 => (x"88",x"c6",x"c1",x"48"),
  1363 => (x"70",x"58",x"a6",x"c4"),
  1364 => (x"e6",x"c0",x"02",x"98"),
  1365 => (x"88",x"c9",x"48",x"87"),
  1366 => (x"70",x"58",x"a6",x"c4"),
  1367 => (x"cd",x"c4",x"02",x"98"),
  1368 => (x"88",x"c1",x"48",x"87"),
  1369 => (x"70",x"58",x"a6",x"c4"),
  1370 => (x"e0",x"c1",x"02",x"98"),
  1371 => (x"88",x"c4",x"48",x"87"),
  1372 => (x"98",x"70",x"58",x"a6"),
  1373 => (x"87",x"f6",x"c3",x"02"),
  1374 => (x"d8",x"87",x"c4",x"c9"),
  1375 => (x"c2",x"c1",x"05",x"66"),
  1376 => (x"48",x"d4",x"ff",x"87"),
  1377 => (x"c0",x"78",x"ff",x"c3"),
  1378 => (x"75",x"1e",x"ca",x"1e"),
  1379 => (x"c1",x"93",x"cb",x"4b"),
  1380 => (x"c4",x"83",x"66",x"c0"),
  1381 => (x"49",x"6c",x"4c",x"a3"),
  1382 => (x"87",x"fe",x"db",x"ff"),
  1383 => (x"1e",x"de",x"1e",x"c1"),
  1384 => (x"db",x"ff",x"49",x"6c"),
  1385 => (x"86",x"d0",x"87",x"f4"),
  1386 => (x"7b",x"c5",x"cc",x"c1"),
  1387 => (x"ad",x"b7",x"66",x"d0"),
  1388 => (x"c1",x"87",x"c5",x"04"),
  1389 => (x"87",x"ce",x"c8",x"85"),
  1390 => (x"c1",x"48",x"66",x"d0"),
  1391 => (x"58",x"a6",x"d4",x"88"),
  1392 => (x"ff",x"87",x"c3",x"c8"),
  1393 => (x"d8",x"87",x"fc",x"da"),
  1394 => (x"f9",x"c7",x"58",x"a6"),
  1395 => (x"c3",x"dd",x"ff",x"87"),
  1396 => (x"58",x"a6",x"cc",x"87"),
  1397 => (x"a8",x"b7",x"66",x"cc"),
  1398 => (x"cc",x"87",x"c6",x"06"),
  1399 => (x"66",x"c8",x"48",x"a6"),
  1400 => (x"ef",x"dc",x"ff",x"78"),
  1401 => (x"a8",x"ec",x"c0",x"87"),
  1402 => (x"87",x"c2",x"c2",x"05"),
  1403 => (x"c1",x"05",x"66",x"d8"),
  1404 => (x"49",x"75",x"87",x"f2"),
  1405 => (x"f8",x"c0",x"91",x"cb"),
  1406 => (x"a1",x"c4",x"81",x"66"),
  1407 => (x"c8",x"4c",x"6a",x"4a"),
  1408 => (x"66",x"c8",x"4a",x"a1"),
  1409 => (x"d3",x"cc",x"c1",x"52"),
  1410 => (x"48",x"d4",x"ff",x"79"),
  1411 => (x"d4",x"78",x"ff",x"c3"),
  1412 => (x"d4",x"ff",x"48",x"a6"),
  1413 => (x"66",x"d4",x"78",x"bf"),
  1414 => (x"87",x"e8",x"c0",x"02"),
  1415 => (x"a8",x"fb",x"c0",x"48"),
  1416 => (x"87",x"e0",x"c0",x"02"),
  1417 => (x"7c",x"97",x"66",x"d4"),
  1418 => (x"d4",x"ff",x"84",x"c1"),
  1419 => (x"78",x"ff",x"c3",x"48"),
  1420 => (x"ff",x"48",x"a6",x"d4"),
  1421 => (x"d4",x"78",x"bf",x"d4"),
  1422 => (x"87",x"c8",x"02",x"66"),
  1423 => (x"a8",x"fb",x"c0",x"48"),
  1424 => (x"87",x"e0",x"ff",x"05"),
  1425 => (x"c2",x"54",x"e0",x"c0"),
  1426 => (x"97",x"c0",x"54",x"c1"),
  1427 => (x"b7",x"66",x"d0",x"7c"),
  1428 => (x"87",x"c5",x"04",x"ad"),
  1429 => (x"ed",x"c5",x"85",x"c1"),
  1430 => (x"48",x"66",x"d0",x"87"),
  1431 => (x"a6",x"d4",x"88",x"c1"),
  1432 => (x"87",x"e2",x"c5",x"58"),
  1433 => (x"87",x"db",x"d8",x"ff"),
  1434 => (x"c5",x"58",x"a6",x"d8"),
  1435 => (x"66",x"c8",x"87",x"d8"),
  1436 => (x"a8",x"66",x"d8",x"48"),
  1437 => (x"87",x"fd",x"c4",x"05"),
  1438 => (x"c0",x"48",x"a6",x"dc"),
  1439 => (x"d3",x"da",x"ff",x"78"),
  1440 => (x"58",x"a6",x"d8",x"87"),
  1441 => (x"87",x"cc",x"da",x"ff"),
  1442 => (x"58",x"a6",x"e4",x"c0"),
  1443 => (x"05",x"a8",x"ec",x"c0"),
  1444 => (x"c0",x"87",x"ca",x"c0"),
  1445 => (x"d4",x"48",x"a6",x"e0"),
  1446 => (x"c6",x"c0",x"78",x"66"),
  1447 => (x"48",x"d4",x"ff",x"87"),
  1448 => (x"75",x"78",x"ff",x"c3"),
  1449 => (x"c0",x"91",x"cb",x"49"),
  1450 => (x"71",x"48",x"66",x"f8"),
  1451 => (x"58",x"a6",x"c4",x"80"),
  1452 => (x"81",x"ca",x"49",x"6e"),
  1453 => (x"c0",x"51",x"66",x"d4"),
  1454 => (x"c1",x"49",x"66",x"e0"),
  1455 => (x"89",x"66",x"d4",x"81"),
  1456 => (x"30",x"71",x"48",x"c1"),
  1457 => (x"89",x"c1",x"49",x"70"),
  1458 => (x"82",x"c8",x"4a",x"6e"),
  1459 => (x"79",x"97",x"09",x"72"),
  1460 => (x"e8",x"e0",x"c2",x"09"),
  1461 => (x"66",x"d4",x"49",x"bf"),
  1462 => (x"6a",x"97",x"29",x"b7"),
  1463 => (x"98",x"71",x"48",x"4a"),
  1464 => (x"58",x"a6",x"e8",x"c0"),
  1465 => (x"80",x"c4",x"48",x"6e"),
  1466 => (x"c4",x"58",x"a6",x"c8"),
  1467 => (x"d8",x"4c",x"bf",x"66"),
  1468 => (x"66",x"c8",x"48",x"66"),
  1469 => (x"c9",x"c0",x"02",x"a8"),
  1470 => (x"a6",x"e0",x"c0",x"87"),
  1471 => (x"c0",x"78",x"c0",x"48"),
  1472 => (x"e0",x"c0",x"87",x"c6"),
  1473 => (x"78",x"c1",x"48",x"a6"),
  1474 => (x"1e",x"66",x"e0",x"c0"),
  1475 => (x"74",x"1e",x"e0",x"c0"),
  1476 => (x"c5",x"d6",x"ff",x"49"),
  1477 => (x"d8",x"86",x"c8",x"87"),
  1478 => (x"b7",x"c0",x"58",x"a6"),
  1479 => (x"da",x"c1",x"06",x"a8"),
  1480 => (x"84",x"66",x"d4",x"87"),
  1481 => (x"49",x"bf",x"66",x"c4"),
  1482 => (x"74",x"81",x"e0",x"c0"),
  1483 => (x"c3",x"c1",x"4b",x"89"),
  1484 => (x"fe",x"71",x"4a",x"c2"),
  1485 => (x"c2",x"87",x"f9",x"e5"),
  1486 => (x"48",x"66",x"dc",x"84"),
  1487 => (x"e0",x"c0",x"80",x"c1"),
  1488 => (x"e4",x"c0",x"58",x"a6"),
  1489 => (x"81",x"c1",x"49",x"66"),
  1490 => (x"c0",x"02",x"a9",x"70"),
  1491 => (x"e0",x"c0",x"87",x"c9"),
  1492 => (x"78",x"c0",x"48",x"a6"),
  1493 => (x"c0",x"87",x"c6",x"c0"),
  1494 => (x"c1",x"48",x"a6",x"e0"),
  1495 => (x"66",x"e0",x"c0",x"78"),
  1496 => (x"bf",x"66",x"c8",x"1e"),
  1497 => (x"81",x"e0",x"c0",x"49"),
  1498 => (x"1e",x"71",x"89",x"74"),
  1499 => (x"d4",x"ff",x"49",x"74"),
  1500 => (x"86",x"c8",x"87",x"e8"),
  1501 => (x"01",x"a8",x"b7",x"c0"),
  1502 => (x"dc",x"87",x"fe",x"fe"),
  1503 => (x"d0",x"c0",x"02",x"66"),
  1504 => (x"c9",x"49",x"6e",x"87"),
  1505 => (x"51",x"66",x"dc",x"81"),
  1506 => (x"cc",x"c1",x"48",x"6e"),
  1507 => (x"cc",x"c0",x"78",x"f4"),
  1508 => (x"c9",x"49",x"6e",x"87"),
  1509 => (x"6e",x"51",x"c2",x"81"),
  1510 => (x"da",x"d0",x"c1",x"48"),
  1511 => (x"b7",x"66",x"d0",x"78"),
  1512 => (x"c5",x"c0",x"04",x"ad"),
  1513 => (x"c0",x"85",x"c1",x"87"),
  1514 => (x"66",x"d0",x"87",x"dc"),
  1515 => (x"d4",x"88",x"c1",x"48"),
  1516 => (x"d1",x"c0",x"58",x"a6"),
  1517 => (x"ca",x"d3",x"ff",x"87"),
  1518 => (x"58",x"a6",x"d8",x"87"),
  1519 => (x"ff",x"87",x"c7",x"c0"),
  1520 => (x"d8",x"87",x"c0",x"d3"),
  1521 => (x"66",x"d4",x"58",x"a6"),
  1522 => (x"87",x"c9",x"c0",x"02"),
  1523 => (x"b7",x"66",x"c0",x"c1"),
  1524 => (x"e4",x"f5",x"04",x"ad"),
  1525 => (x"ad",x"b7",x"c7",x"87"),
  1526 => (x"87",x"d9",x"c0",x"03"),
  1527 => (x"91",x"cb",x"49",x"75"),
  1528 => (x"81",x"66",x"f8",x"c0"),
  1529 => (x"6a",x"4a",x"a1",x"c4"),
  1530 => (x"79",x"52",x"c0",x"4a"),
  1531 => (x"b7",x"c7",x"85",x"c1"),
  1532 => (x"e7",x"ff",x"04",x"ad"),
  1533 => (x"02",x"66",x"d8",x"87"),
  1534 => (x"c0",x"87",x"e2",x"c0"),
  1535 => (x"c1",x"49",x"66",x"f8"),
  1536 => (x"f8",x"c0",x"81",x"cd"),
  1537 => (x"d5",x"c1",x"4a",x"66"),
  1538 => (x"c1",x"52",x"c0",x"82"),
  1539 => (x"c0",x"79",x"d3",x"cc"),
  1540 => (x"c1",x"49",x"66",x"f8"),
  1541 => (x"c3",x"c1",x"81",x"d1"),
  1542 => (x"d6",x"c0",x"79",x"c5"),
  1543 => (x"66",x"f8",x"c0",x"87"),
  1544 => (x"81",x"cd",x"c1",x"49"),
  1545 => (x"4a",x"66",x"f8",x"c0"),
  1546 => (x"c1",x"82",x"d1",x"c1"),
  1547 => (x"c2",x"7a",x"cc",x"c3"),
  1548 => (x"c1",x"79",x"f2",x"c8"),
  1549 => (x"c0",x"4a",x"eb",x"d0"),
  1550 => (x"c1",x"49",x"66",x"f8"),
  1551 => (x"79",x"72",x"81",x"d8"),
  1552 => (x"48",x"bf",x"d0",x"ff"),
  1553 => (x"98",x"c0",x"c0",x"c8"),
  1554 => (x"70",x"58",x"a6",x"c4"),
  1555 => (x"d1",x"c0",x"02",x"98"),
  1556 => (x"bf",x"d0",x"ff",x"87"),
  1557 => (x"c0",x"c0",x"c8",x"48"),
  1558 => (x"58",x"a6",x"c4",x"98"),
  1559 => (x"ff",x"05",x"98",x"70"),
  1560 => (x"d0",x"ff",x"87",x"ef"),
  1561 => (x"78",x"e0",x"c0",x"48"),
  1562 => (x"ff",x"48",x"66",x"cc"),
  1563 => (x"d2",x"ff",x"8e",x"d8"),
  1564 => (x"c7",x"1e",x"87",x"da"),
  1565 => (x"c1",x"1e",x"c0",x"1e"),
  1566 => (x"c2",x"1e",x"f8",x"e3"),
  1567 => (x"49",x"bf",x"ec",x"e0"),
  1568 => (x"c1",x"87",x"ed",x"ef"),
  1569 => (x"c0",x"49",x"f8",x"e3"),
  1570 => (x"f4",x"87",x"d4",x"e6"),
  1571 => (x"1e",x"4f",x"26",x"8e"),
  1572 => (x"c2",x"87",x"fd",x"c9"),
  1573 => (x"c0",x"48",x"c8",x"e1"),
  1574 => (x"48",x"d4",x"ff",x"50"),
  1575 => (x"c1",x"78",x"ff",x"c3"),
  1576 => (x"fe",x"49",x"d3",x"c3"),
  1577 => (x"fe",x"87",x"e5",x"df"),
  1578 => (x"70",x"87",x"f0",x"e8"),
  1579 => (x"87",x"cd",x"02",x"98"),
  1580 => (x"87",x"ed",x"f4",x"fe"),
  1581 => (x"c4",x"02",x"98",x"70"),
  1582 => (x"c2",x"4a",x"c1",x"87"),
  1583 => (x"72",x"4a",x"c0",x"87"),
  1584 => (x"87",x"c8",x"02",x"9a"),
  1585 => (x"49",x"dd",x"c3",x"c1"),
  1586 => (x"87",x"c0",x"df",x"fe"),
  1587 => (x"bf",x"f4",x"e3",x"c1"),
  1588 => (x"cb",x"d6",x"ff",x"49"),
  1589 => (x"c0",x"e1",x"c2",x"87"),
  1590 => (x"c2",x"78",x"c0",x"48"),
  1591 => (x"c0",x"48",x"ec",x"e0"),
  1592 => (x"cd",x"fe",x"49",x"78"),
  1593 => (x"87",x"d4",x"c3",x"87"),
  1594 => (x"c0",x"87",x"f9",x"c8"),
  1595 => (x"ff",x"87",x"d2",x"e5"),
  1596 => (x"4f",x"26",x"87",x"f6"),
  1597 => (x"00",x"00",x"10",x"e0"),
  1598 => (x"00",x"00",x"10",x"42"),
  1599 => (x"00",x"00",x"28",x"58"),
  1600 => (x"42",x"00",x"00",x"00"),
  1601 => (x"76",x"00",x"00",x"10"),
  1602 => (x"00",x"00",x"00",x"28"),
  1603 => (x"10",x"42",x"00",x"00"),
  1604 => (x"28",x"94",x"00",x"00"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"10",x"42",x"00"),
  1607 => (x"00",x"28",x"b2",x"00"),
  1608 => (x"00",x"00",x"00",x"00"),
  1609 => (x"00",x"00",x"10",x"42"),
  1610 => (x"00",x"00",x"28",x"d0"),
  1611 => (x"42",x"00",x"00",x"00"),
  1612 => (x"ee",x"00",x"00",x"10"),
  1613 => (x"00",x"00",x"00",x"28"),
  1614 => (x"10",x"42",x"00",x"00"),
  1615 => (x"29",x"0c",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"13",x"13",x"00"),
  1618 => (x"00",x"00",x"00",x"00"),
  1619 => (x"00",x"00",x"00",x"00"),
  1620 => (x"00",x"00",x"11",x"12"),
  1621 => (x"00",x"00",x"00",x"00"),
  1622 => (x"1e",x"00",x"00",x"00"),
  1623 => (x"87",x"d5",x"c1",x"1e"),
  1624 => (x"26",x"58",x"a6",x"c4"),
  1625 => (x"71",x"1e",x"4f",x"26"),
  1626 => (x"48",x"f0",x"fe",x"4a"),
  1627 => (x"0a",x"cd",x"78",x"c0"),
  1628 => (x"e5",x"c1",x"0a",x"7a"),
  1629 => (x"dc",x"fe",x"49",x"fc"),
  1630 => (x"4f",x"26",x"87",x"d2"),
  1631 => (x"20",x"74",x"65",x"53"),
  1632 => (x"64",x"6e",x"61",x"68"),
  1633 => (x"0a",x"72",x"65",x"6c"),
  1634 => (x"20",x"6e",x"49",x"00"),
  1635 => (x"65",x"74",x"6e",x"69"),
  1636 => (x"70",x"75",x"72",x"72"),
  1637 => (x"6f",x"63",x"20",x"74"),
  1638 => (x"72",x"74",x"73",x"6e"),
  1639 => (x"6f",x"74",x"63",x"75"),
  1640 => (x"1e",x"00",x"0a",x"72"),
  1641 => (x"49",x"c9",x"e6",x"c1"),
  1642 => (x"87",x"e0",x"db",x"fe"),
  1643 => (x"49",x"db",x"e5",x"c1"),
  1644 => (x"26",x"87",x"f3",x"fe"),
  1645 => (x"f0",x"fe",x"1e",x"4f"),
  1646 => (x"4f",x"26",x"48",x"bf"),
  1647 => (x"48",x"f0",x"fe",x"1e"),
  1648 => (x"4f",x"26",x"78",x"c1"),
  1649 => (x"48",x"f0",x"fe",x"1e"),
  1650 => (x"4f",x"26",x"78",x"c0"),
  1651 => (x"c0",x"4a",x"71",x"1e"),
  1652 => (x"49",x"a2",x"c4",x"7a"),
  1653 => (x"a2",x"c8",x"79",x"c0"),
  1654 => (x"cc",x"79",x"c0",x"49"),
  1655 => (x"79",x"c0",x"49",x"a2"),
  1656 => (x"5e",x"0e",x"4f",x"26"),
  1657 => (x"f8",x"0e",x"5c",x"5b"),
  1658 => (x"c8",x"4c",x"71",x"86"),
  1659 => (x"a4",x"cc",x"49",x"a4"),
  1660 => (x"c1",x"48",x"6b",x"4b"),
  1661 => (x"58",x"a6",x"c4",x"80"),
  1662 => (x"a6",x"c8",x"98",x"cf"),
  1663 => (x"c4",x"48",x"69",x"58"),
  1664 => (x"d4",x"05",x"a8",x"66"),
  1665 => (x"c1",x"48",x"6b",x"87"),
  1666 => (x"58",x"a6",x"c4",x"80"),
  1667 => (x"a6",x"c8",x"98",x"cf"),
  1668 => (x"c4",x"48",x"69",x"58"),
  1669 => (x"ec",x"02",x"a8",x"66"),
  1670 => (x"87",x"e8",x"fe",x"87"),
  1671 => (x"49",x"a4",x"d0",x"c1"),
  1672 => (x"90",x"c4",x"48",x"6b"),
  1673 => (x"70",x"58",x"a6",x"c4"),
  1674 => (x"79",x"66",x"d4",x"81"),
  1675 => (x"80",x"c1",x"48",x"6b"),
  1676 => (x"cf",x"58",x"a6",x"c8"),
  1677 => (x"c1",x"7b",x"70",x"98"),
  1678 => (x"ff",x"fd",x"87",x"d2"),
  1679 => (x"c2",x"8e",x"f8",x"87"),
  1680 => (x"26",x"4d",x"26",x"87"),
  1681 => (x"26",x"4b",x"26",x"4c"),
  1682 => (x"5b",x"5e",x"0e",x"4f"),
  1683 => (x"f8",x"0e",x"5d",x"5c"),
  1684 => (x"c4",x"4d",x"71",x"86"),
  1685 => (x"48",x"6d",x"4c",x"a5"),
  1686 => (x"c5",x"05",x"a8",x"6c"),
  1687 => (x"c0",x"48",x"ff",x"87"),
  1688 => (x"df",x"fd",x"87",x"e5"),
  1689 => (x"4b",x"a5",x"d0",x"87"),
  1690 => (x"90",x"c4",x"48",x"6c"),
  1691 => (x"70",x"58",x"a6",x"c4"),
  1692 => (x"c3",x"4b",x"6b",x"83"),
  1693 => (x"48",x"6c",x"9b",x"ff"),
  1694 => (x"a6",x"c8",x"80",x"c1"),
  1695 => (x"70",x"98",x"cf",x"58"),
  1696 => (x"87",x"f8",x"fc",x"7c"),
  1697 => (x"f8",x"48",x"49",x"73"),
  1698 => (x"87",x"f5",x"fe",x"8e"),
  1699 => (x"f8",x"1e",x"73",x"1e"),
  1700 => (x"87",x"f0",x"fc",x"86"),
  1701 => (x"49",x"4b",x"bf",x"e0"),
  1702 => (x"99",x"c0",x"e0",x"c0"),
  1703 => (x"87",x"e7",x"c0",x"02"),
  1704 => (x"ff",x"c3",x"4a",x"73"),
  1705 => (x"ea",x"e4",x"c2",x"9a"),
  1706 => (x"90",x"c4",x"48",x"bf"),
  1707 => (x"c2",x"58",x"a6",x"c4"),
  1708 => (x"70",x"49",x"fa",x"e4"),
  1709 => (x"c2",x"79",x"72",x"81"),
  1710 => (x"48",x"bf",x"ea",x"e4"),
  1711 => (x"a6",x"c8",x"80",x"c1"),
  1712 => (x"c2",x"98",x"cf",x"58"),
  1713 => (x"73",x"58",x"ee",x"e4"),
  1714 => (x"99",x"c0",x"d0",x"49"),
  1715 => (x"87",x"f2",x"c0",x"02"),
  1716 => (x"bf",x"f2",x"e4",x"c2"),
  1717 => (x"f6",x"e4",x"c2",x"48"),
  1718 => (x"c0",x"02",x"a8",x"bf"),
  1719 => (x"e4",x"c2",x"87",x"e4"),
  1720 => (x"c4",x"48",x"bf",x"f2"),
  1721 => (x"58",x"a6",x"c4",x"90"),
  1722 => (x"49",x"fa",x"e5",x"c2"),
  1723 => (x"48",x"e0",x"81",x"70"),
  1724 => (x"e4",x"c2",x"78",x"69"),
  1725 => (x"c1",x"48",x"bf",x"f2"),
  1726 => (x"58",x"a6",x"c8",x"80"),
  1727 => (x"e4",x"c2",x"98",x"cf"),
  1728 => (x"f0",x"fa",x"58",x"f6"),
  1729 => (x"58",x"a6",x"c4",x"87"),
  1730 => (x"f8",x"87",x"f1",x"fa"),
  1731 => (x"87",x"f5",x"fc",x"8e"),
  1732 => (x"ea",x"e4",x"c2",x"1e"),
  1733 => (x"87",x"f4",x"fa",x"49"),
  1734 => (x"49",x"cc",x"ea",x"c1"),
  1735 => (x"c3",x"87",x"c7",x"f9"),
  1736 => (x"4f",x"26",x"87",x"f5"),
  1737 => (x"c2",x"1e",x"73",x"1e"),
  1738 => (x"fc",x"49",x"ea",x"e4"),
  1739 => (x"4a",x"70",x"87",x"db"),
  1740 => (x"04",x"aa",x"b7",x"c0"),
  1741 => (x"c3",x"87",x"cc",x"c2"),
  1742 => (x"c9",x"05",x"aa",x"f0"),
  1743 => (x"cf",x"ef",x"c1",x"87"),
  1744 => (x"c1",x"78",x"c1",x"48"),
  1745 => (x"e0",x"c3",x"87",x"ed"),
  1746 => (x"87",x"c9",x"05",x"aa"),
  1747 => (x"48",x"d3",x"ef",x"c1"),
  1748 => (x"de",x"c1",x"78",x"c1"),
  1749 => (x"d3",x"ef",x"c1",x"87"),
  1750 => (x"87",x"c6",x"02",x"bf"),
  1751 => (x"4b",x"a2",x"c0",x"c2"),
  1752 => (x"4b",x"72",x"87",x"c2"),
  1753 => (x"bf",x"cf",x"ef",x"c1"),
  1754 => (x"87",x"e0",x"c0",x"02"),
  1755 => (x"b7",x"c4",x"49",x"73"),
  1756 => (x"ef",x"c1",x"91",x"29"),
  1757 => (x"4a",x"73",x"81",x"d7"),
  1758 => (x"92",x"c2",x"9a",x"cf"),
  1759 => (x"30",x"72",x"48",x"c1"),
  1760 => (x"ba",x"ff",x"4a",x"70"),
  1761 => (x"98",x"69",x"48",x"72"),
  1762 => (x"87",x"db",x"79",x"70"),
  1763 => (x"b7",x"c4",x"49",x"73"),
  1764 => (x"ef",x"c1",x"91",x"29"),
  1765 => (x"4a",x"73",x"81",x"d7"),
  1766 => (x"92",x"c2",x"9a",x"cf"),
  1767 => (x"30",x"72",x"48",x"c3"),
  1768 => (x"69",x"48",x"4a",x"70"),
  1769 => (x"c1",x"79",x"70",x"b0"),
  1770 => (x"c0",x"48",x"d3",x"ef"),
  1771 => (x"cf",x"ef",x"c1",x"78"),
  1772 => (x"c2",x"78",x"c0",x"48"),
  1773 => (x"fa",x"49",x"ea",x"e4"),
  1774 => (x"4a",x"70",x"87",x"cf"),
  1775 => (x"03",x"aa",x"b7",x"c0"),
  1776 => (x"c0",x"87",x"f4",x"fd"),
  1777 => (x"26",x"87",x"c4",x"48"),
  1778 => (x"26",x"4c",x"26",x"4d"),
  1779 => (x"00",x"4f",x"26",x"4b"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"1e",x"00",x"00",x"00"),
  1798 => (x"49",x"72",x"4a",x"c0"),
  1799 => (x"ef",x"c1",x"91",x"c4"),
  1800 => (x"79",x"c0",x"81",x"d7"),
  1801 => (x"b7",x"d0",x"82",x"c1"),
  1802 => (x"87",x"ee",x"04",x"aa"),
  1803 => (x"5e",x"0e",x"4f",x"26"),
  1804 => (x"0e",x"5d",x"5c",x"5b"),
  1805 => (x"cb",x"f6",x"4d",x"71"),
  1806 => (x"c4",x"4a",x"75",x"87"),
  1807 => (x"c1",x"92",x"2a",x"b7"),
  1808 => (x"75",x"82",x"d7",x"ef"),
  1809 => (x"c2",x"9c",x"cf",x"4c"),
  1810 => (x"4b",x"49",x"6a",x"94"),
  1811 => (x"9b",x"c3",x"2b",x"74"),
  1812 => (x"30",x"74",x"48",x"c2"),
  1813 => (x"bc",x"ff",x"4c",x"70"),
  1814 => (x"98",x"71",x"48",x"74"),
  1815 => (x"db",x"f5",x"7a",x"70"),
  1816 => (x"fd",x"48",x"73",x"87"),
  1817 => (x"1e",x"1e",x"87",x"e1"),
  1818 => (x"48",x"bf",x"d0",x"ff"),
  1819 => (x"98",x"c0",x"c0",x"c8"),
  1820 => (x"70",x"58",x"a6",x"c4"),
  1821 => (x"87",x"d0",x"02",x"98"),
  1822 => (x"48",x"bf",x"d0",x"ff"),
  1823 => (x"98",x"c0",x"c0",x"c8"),
  1824 => (x"70",x"58",x"a6",x"c4"),
  1825 => (x"87",x"f0",x"05",x"98"),
  1826 => (x"c4",x"48",x"d0",x"ff"),
  1827 => (x"48",x"71",x"78",x"e1"),
  1828 => (x"78",x"08",x"d4",x"ff"),
  1829 => (x"ff",x"48",x"66",x"c8"),
  1830 => (x"26",x"78",x"08",x"d4"),
  1831 => (x"1e",x"1e",x"4f",x"26"),
  1832 => (x"66",x"c8",x"4a",x"71"),
  1833 => (x"49",x"72",x"1e",x"49"),
  1834 => (x"c4",x"87",x"fb",x"fe"),
  1835 => (x"bf",x"d0",x"ff",x"86"),
  1836 => (x"c0",x"c0",x"c8",x"48"),
  1837 => (x"58",x"a6",x"c4",x"98"),
  1838 => (x"d0",x"02",x"98",x"70"),
  1839 => (x"bf",x"d0",x"ff",x"87"),
  1840 => (x"c0",x"c0",x"c8",x"48"),
  1841 => (x"58",x"a6",x"c4",x"98"),
  1842 => (x"f0",x"05",x"98",x"70"),
  1843 => (x"48",x"d0",x"ff",x"87"),
  1844 => (x"26",x"78",x"e0",x"c0"),
  1845 => (x"73",x"1e",x"4f",x"26"),
  1846 => (x"c8",x"4b",x"71",x"1e"),
  1847 => (x"4a",x"73",x"1e",x"66"),
  1848 => (x"49",x"a2",x"e0",x"c1"),
  1849 => (x"26",x"87",x"f7",x"fe"),
  1850 => (x"4d",x"26",x"87",x"c4"),
  1851 => (x"4b",x"26",x"4c",x"26"),
  1852 => (x"1e",x"1e",x"4f",x"26"),
  1853 => (x"48",x"bf",x"d0",x"ff"),
  1854 => (x"98",x"c0",x"c0",x"c8"),
  1855 => (x"70",x"58",x"a6",x"c4"),
  1856 => (x"87",x"d0",x"02",x"98"),
  1857 => (x"48",x"bf",x"d0",x"ff"),
  1858 => (x"98",x"c0",x"c0",x"c8"),
  1859 => (x"70",x"58",x"a6",x"c4"),
  1860 => (x"87",x"f0",x"05",x"98"),
  1861 => (x"c4",x"48",x"d0",x"ff"),
  1862 => (x"48",x"71",x"78",x"c9"),
  1863 => (x"78",x"08",x"d4",x"ff"),
  1864 => (x"1e",x"4f",x"26",x"26"),
  1865 => (x"49",x"4a",x"71",x"1e"),
  1866 => (x"ff",x"87",x"c7",x"ff"),
  1867 => (x"c8",x"48",x"bf",x"d0"),
  1868 => (x"c4",x"98",x"c0",x"c0"),
  1869 => (x"98",x"70",x"58",x"a6"),
  1870 => (x"ff",x"87",x"d0",x"02"),
  1871 => (x"c8",x"48",x"bf",x"d0"),
  1872 => (x"c4",x"98",x"c0",x"c0"),
  1873 => (x"98",x"70",x"58",x"a6"),
  1874 => (x"ff",x"87",x"f0",x"05"),
  1875 => (x"78",x"c8",x"48",x"d0"),
  1876 => (x"1e",x"4f",x"26",x"26"),
  1877 => (x"71",x"1e",x"1e",x"73"),
  1878 => (x"c6",x"e7",x"c2",x"4b"),
  1879 => (x"87",x"c3",x"02",x"bf"),
  1880 => (x"ff",x"87",x"cc",x"c3"),
  1881 => (x"c8",x"48",x"bf",x"d0"),
  1882 => (x"c4",x"98",x"c0",x"c0"),
  1883 => (x"98",x"70",x"58",x"a6"),
  1884 => (x"ff",x"87",x"d0",x"02"),
  1885 => (x"c8",x"48",x"bf",x"d0"),
  1886 => (x"c4",x"98",x"c0",x"c0"),
  1887 => (x"98",x"70",x"58",x"a6"),
  1888 => (x"ff",x"87",x"f0",x"05"),
  1889 => (x"c9",x"c4",x"48",x"d0"),
  1890 => (x"c0",x"48",x"73",x"78"),
  1891 => (x"d4",x"ff",x"b0",x"e0"),
  1892 => (x"e6",x"c2",x"78",x"08"),
  1893 => (x"78",x"c0",x"48",x"fa"),
  1894 => (x"c5",x"02",x"66",x"cc"),
  1895 => (x"49",x"ff",x"c3",x"87"),
  1896 => (x"49",x"c0",x"87",x"c2"),
  1897 => (x"59",x"c2",x"e7",x"c2"),
  1898 => (x"c6",x"02",x"66",x"d0"),
  1899 => (x"d5",x"d5",x"c5",x"87"),
  1900 => (x"cf",x"87",x"c4",x"4a"),
  1901 => (x"c2",x"4a",x"ff",x"ff"),
  1902 => (x"c2",x"5a",x"c6",x"e7"),
  1903 => (x"c1",x"48",x"c6",x"e7"),
  1904 => (x"87",x"c4",x"26",x"78"),
  1905 => (x"4c",x"26",x"4d",x"26"),
  1906 => (x"4f",x"26",x"4b",x"26"),
  1907 => (x"5c",x"5b",x"5e",x"0e"),
  1908 => (x"4a",x"71",x"0e",x"5d"),
  1909 => (x"bf",x"c2",x"e7",x"c2"),
  1910 => (x"02",x"9a",x"72",x"4c"),
  1911 => (x"c8",x"49",x"87",x"cb"),
  1912 => (x"cd",x"f6",x"c1",x"91"),
  1913 => (x"c4",x"83",x"71",x"4b"),
  1914 => (x"cd",x"fa",x"c1",x"87"),
  1915 => (x"13",x"4d",x"c0",x"4b"),
  1916 => (x"c2",x"99",x"74",x"49"),
  1917 => (x"48",x"bf",x"fe",x"e6"),
  1918 => (x"d4",x"ff",x"b8",x"71"),
  1919 => (x"b7",x"c1",x"78",x"08"),
  1920 => (x"b7",x"c8",x"85",x"2c"),
  1921 => (x"87",x"e7",x"04",x"ad"),
  1922 => (x"bf",x"fa",x"e6",x"c2"),
  1923 => (x"c2",x"80",x"c8",x"48"),
  1924 => (x"fe",x"58",x"fe",x"e6"),
  1925 => (x"73",x"1e",x"87",x"ee"),
  1926 => (x"13",x"4b",x"71",x"1e"),
  1927 => (x"cb",x"02",x"9a",x"4a"),
  1928 => (x"fe",x"49",x"72",x"87"),
  1929 => (x"4a",x"13",x"87",x"e6"),
  1930 => (x"87",x"f5",x"05",x"9a"),
  1931 => (x"1e",x"87",x"d9",x"fe"),
  1932 => (x"fa",x"e6",x"c2",x"1e"),
  1933 => (x"e6",x"c2",x"49",x"bf"),
  1934 => (x"a1",x"c1",x"48",x"fa"),
  1935 => (x"b7",x"c0",x"c4",x"78"),
  1936 => (x"87",x"db",x"03",x"a9"),
  1937 => (x"c2",x"48",x"d4",x"ff"),
  1938 => (x"78",x"bf",x"fe",x"e6"),
  1939 => (x"bf",x"fa",x"e6",x"c2"),
  1940 => (x"fa",x"e6",x"c2",x"49"),
  1941 => (x"78",x"a1",x"c1",x"48"),
  1942 => (x"a9",x"b7",x"c0",x"c4"),
  1943 => (x"ff",x"87",x"e5",x"04"),
  1944 => (x"c8",x"48",x"bf",x"d0"),
  1945 => (x"c4",x"98",x"c0",x"c0"),
  1946 => (x"98",x"70",x"58",x"a6"),
  1947 => (x"ff",x"87",x"d0",x"02"),
  1948 => (x"c8",x"48",x"bf",x"d0"),
  1949 => (x"c4",x"98",x"c0",x"c0"),
  1950 => (x"98",x"70",x"58",x"a6"),
  1951 => (x"ff",x"87",x"f0",x"05"),
  1952 => (x"78",x"c8",x"48",x"d0"),
  1953 => (x"48",x"c6",x"e7",x"c2"),
  1954 => (x"26",x"26",x"78",x"c0"),
  1955 => (x"00",x"00",x"00",x"4f"),
  1956 => (x"00",x"00",x"00",x"00"),
  1957 => (x"00",x"00",x"00",x"00"),
  1958 => (x"00",x"00",x"5f",x"5f"),
  1959 => (x"03",x"03",x"00",x"00"),
  1960 => (x"00",x"03",x"03",x"00"),
  1961 => (x"7f",x"7f",x"14",x"00"),
  1962 => (x"14",x"7f",x"7f",x"14"),
  1963 => (x"2e",x"24",x"00",x"00"),
  1964 => (x"12",x"3a",x"6b",x"6b"),
  1965 => (x"36",x"6a",x"4c",x"00"),
  1966 => (x"32",x"56",x"6c",x"18"),
  1967 => (x"4f",x"7e",x"30",x"00"),
  1968 => (x"68",x"3a",x"77",x"59"),
  1969 => (x"04",x"00",x"00",x"40"),
  1970 => (x"00",x"00",x"03",x"07"),
  1971 => (x"1c",x"00",x"00",x"00"),
  1972 => (x"00",x"41",x"63",x"3e"),
  1973 => (x"41",x"00",x"00",x"00"),
  1974 => (x"00",x"1c",x"3e",x"63"),
  1975 => (x"3e",x"2a",x"08",x"00"),
  1976 => (x"2a",x"3e",x"1c",x"1c"),
  1977 => (x"08",x"08",x"00",x"08"),
  1978 => (x"08",x"08",x"3e",x"3e"),
  1979 => (x"80",x"00",x"00",x"00"),
  1980 => (x"00",x"00",x"60",x"e0"),
  1981 => (x"08",x"08",x"00",x"00"),
  1982 => (x"08",x"08",x"08",x"08"),
  1983 => (x"00",x"00",x"00",x"00"),
  1984 => (x"00",x"00",x"60",x"60"),
  1985 => (x"30",x"60",x"40",x"00"),
  1986 => (x"03",x"06",x"0c",x"18"),
  1987 => (x"7f",x"3e",x"00",x"01"),
  1988 => (x"3e",x"7f",x"4d",x"59"),
  1989 => (x"06",x"04",x"00",x"00"),
  1990 => (x"00",x"00",x"7f",x"7f"),
  1991 => (x"63",x"42",x"00",x"00"),
  1992 => (x"46",x"4f",x"59",x"71"),
  1993 => (x"63",x"22",x"00",x"00"),
  1994 => (x"36",x"7f",x"49",x"49"),
  1995 => (x"16",x"1c",x"18",x"00"),
  1996 => (x"10",x"7f",x"7f",x"13"),
  1997 => (x"67",x"27",x"00",x"00"),
  1998 => (x"39",x"7d",x"45",x"45"),
  1999 => (x"7e",x"3c",x"00",x"00"),
  2000 => (x"30",x"79",x"49",x"4b"),
  2001 => (x"01",x"01",x"00",x"00"),
  2002 => (x"07",x"0f",x"79",x"71"),
  2003 => (x"7f",x"36",x"00",x"00"),
  2004 => (x"36",x"7f",x"49",x"49"),
  2005 => (x"4f",x"06",x"00",x"00"),
  2006 => (x"1e",x"3f",x"69",x"49"),
  2007 => (x"00",x"00",x"00",x"00"),
  2008 => (x"00",x"00",x"66",x"66"),
  2009 => (x"80",x"00",x"00",x"00"),
  2010 => (x"00",x"00",x"66",x"e6"),
  2011 => (x"08",x"08",x"00",x"00"),
  2012 => (x"22",x"22",x"14",x"14"),
  2013 => (x"14",x"14",x"00",x"00"),
  2014 => (x"14",x"14",x"14",x"14"),
  2015 => (x"22",x"22",x"00",x"00"),
  2016 => (x"08",x"08",x"14",x"14"),
  2017 => (x"03",x"02",x"00",x"00"),
  2018 => (x"06",x"0f",x"59",x"51"),
  2019 => (x"41",x"7f",x"3e",x"00"),
  2020 => (x"1e",x"1f",x"55",x"5d"),
  2021 => (x"7f",x"7e",x"00",x"00"),
  2022 => (x"7e",x"7f",x"09",x"09"),
  2023 => (x"7f",x"7f",x"00",x"00"),
  2024 => (x"36",x"7f",x"49",x"49"),
  2025 => (x"3e",x"1c",x"00",x"00"),
  2026 => (x"41",x"41",x"41",x"63"),
  2027 => (x"7f",x"7f",x"00",x"00"),
  2028 => (x"1c",x"3e",x"63",x"41"),
  2029 => (x"7f",x"7f",x"00",x"00"),
  2030 => (x"41",x"41",x"49",x"49"),
  2031 => (x"7f",x"7f",x"00",x"00"),
  2032 => (x"01",x"01",x"09",x"09"),
  2033 => (x"7f",x"3e",x"00",x"00"),
  2034 => (x"7a",x"7b",x"49",x"41"),
  2035 => (x"7f",x"7f",x"00",x"00"),
  2036 => (x"7f",x"7f",x"08",x"08"),
  2037 => (x"41",x"00",x"00",x"00"),
  2038 => (x"00",x"41",x"7f",x"7f"),
  2039 => (x"60",x"20",x"00",x"00"),
  2040 => (x"3f",x"7f",x"40",x"40"),
  2041 => (x"08",x"7f",x"7f",x"00"),
  2042 => (x"41",x"63",x"36",x"1c"),
  2043 => (x"7f",x"7f",x"00",x"00"),
  2044 => (x"40",x"40",x"40",x"40"),
  2045 => (x"06",x"7f",x"7f",x"00"),
  2046 => (x"7f",x"7f",x"06",x"0c"),
  2047 => (x"06",x"7f",x"7f",x"00"),
  2048 => (x"7f",x"7f",x"18",x"0c"),
  2049 => (x"7f",x"3e",x"00",x"00"),
  2050 => (x"3e",x"7f",x"41",x"41"),
  2051 => (x"7f",x"7f",x"00",x"00"),
  2052 => (x"06",x"0f",x"09",x"09"),
  2053 => (x"41",x"7f",x"3e",x"00"),
  2054 => (x"40",x"7e",x"7f",x"61"),
  2055 => (x"7f",x"7f",x"00",x"00"),
  2056 => (x"66",x"7f",x"19",x"09"),
  2057 => (x"6f",x"26",x"00",x"00"),
  2058 => (x"32",x"7b",x"59",x"4d"),
  2059 => (x"01",x"01",x"00",x"00"),
  2060 => (x"01",x"01",x"7f",x"7f"),
  2061 => (x"7f",x"3f",x"00",x"00"),
  2062 => (x"3f",x"7f",x"40",x"40"),
  2063 => (x"3f",x"0f",x"00",x"00"),
  2064 => (x"0f",x"3f",x"70",x"70"),
  2065 => (x"30",x"7f",x"7f",x"00"),
  2066 => (x"7f",x"7f",x"30",x"18"),
  2067 => (x"36",x"63",x"41",x"00"),
  2068 => (x"63",x"36",x"1c",x"1c"),
  2069 => (x"06",x"03",x"01",x"41"),
  2070 => (x"03",x"06",x"7c",x"7c"),
  2071 => (x"59",x"71",x"61",x"01"),
  2072 => (x"41",x"43",x"47",x"4d"),
  2073 => (x"7f",x"00",x"00",x"00"),
  2074 => (x"00",x"41",x"41",x"7f"),
  2075 => (x"06",x"03",x"01",x"00"),
  2076 => (x"60",x"30",x"18",x"0c"),
  2077 => (x"41",x"00",x"00",x"40"),
  2078 => (x"00",x"7f",x"7f",x"41"),
  2079 => (x"06",x"0c",x"08",x"00"),
  2080 => (x"08",x"0c",x"06",x"03"),
  2081 => (x"80",x"80",x"80",x"00"),
  2082 => (x"80",x"80",x"80",x"80"),
  2083 => (x"00",x"00",x"00",x"00"),
  2084 => (x"00",x"04",x"07",x"03"),
  2085 => (x"74",x"20",x"00",x"00"),
  2086 => (x"78",x"7c",x"54",x"54"),
  2087 => (x"7f",x"7f",x"00",x"00"),
  2088 => (x"38",x"7c",x"44",x"44"),
  2089 => (x"7c",x"38",x"00",x"00"),
  2090 => (x"00",x"44",x"44",x"44"),
  2091 => (x"7c",x"38",x"00",x"00"),
  2092 => (x"7f",x"7f",x"44",x"44"),
  2093 => (x"7c",x"38",x"00",x"00"),
  2094 => (x"18",x"5c",x"54",x"54"),
  2095 => (x"7e",x"04",x"00",x"00"),
  2096 => (x"00",x"05",x"05",x"7f"),
  2097 => (x"bc",x"18",x"00",x"00"),
  2098 => (x"7c",x"fc",x"a4",x"a4"),
  2099 => (x"7f",x"7f",x"00",x"00"),
  2100 => (x"78",x"7c",x"04",x"04"),
  2101 => (x"00",x"00",x"00",x"00"),
  2102 => (x"00",x"40",x"7d",x"3d"),
  2103 => (x"80",x"80",x"00",x"00"),
  2104 => (x"00",x"7d",x"fd",x"80"),
  2105 => (x"7f",x"7f",x"00",x"00"),
  2106 => (x"44",x"6c",x"38",x"10"),
  2107 => (x"00",x"00",x"00",x"00"),
  2108 => (x"00",x"40",x"7f",x"3f"),
  2109 => (x"0c",x"7c",x"7c",x"00"),
  2110 => (x"78",x"7c",x"0c",x"18"),
  2111 => (x"7c",x"7c",x"00",x"00"),
  2112 => (x"78",x"7c",x"04",x"04"),
  2113 => (x"7c",x"38",x"00",x"00"),
  2114 => (x"38",x"7c",x"44",x"44"),
  2115 => (x"fc",x"fc",x"00",x"00"),
  2116 => (x"18",x"3c",x"24",x"24"),
  2117 => (x"3c",x"18",x"00",x"00"),
  2118 => (x"fc",x"fc",x"24",x"24"),
  2119 => (x"7c",x"7c",x"00",x"00"),
  2120 => (x"08",x"0c",x"04",x"04"),
  2121 => (x"5c",x"48",x"00",x"00"),
  2122 => (x"20",x"74",x"54",x"54"),
  2123 => (x"3f",x"04",x"00",x"00"),
  2124 => (x"00",x"44",x"44",x"7f"),
  2125 => (x"7c",x"3c",x"00",x"00"),
  2126 => (x"7c",x"7c",x"40",x"40"),
  2127 => (x"3c",x"1c",x"00",x"00"),
  2128 => (x"1c",x"3c",x"60",x"60"),
  2129 => (x"60",x"7c",x"3c",x"00"),
  2130 => (x"3c",x"7c",x"60",x"30"),
  2131 => (x"38",x"6c",x"44",x"00"),
  2132 => (x"44",x"6c",x"38",x"10"),
  2133 => (x"bc",x"1c",x"00",x"00"),
  2134 => (x"1c",x"3c",x"60",x"e0"),
  2135 => (x"64",x"44",x"00",x"00"),
  2136 => (x"44",x"4c",x"5c",x"74"),
  2137 => (x"08",x"08",x"00",x"00"),
  2138 => (x"41",x"41",x"77",x"3e"),
  2139 => (x"00",x"00",x"00",x"00"),
  2140 => (x"00",x"00",x"7f",x"7f"),
  2141 => (x"41",x"41",x"00",x"00"),
  2142 => (x"08",x"08",x"3e",x"77"),
  2143 => (x"01",x"01",x"02",x"00"),
  2144 => (x"01",x"02",x"02",x"03"),
  2145 => (x"7f",x"7f",x"7f",x"00"),
  2146 => (x"7f",x"7f",x"7f",x"7f"),
  2147 => (x"1c",x"08",x"08",x"00"),
  2148 => (x"7f",x"3e",x"3e",x"1c"),
  2149 => (x"3e",x"7f",x"7f",x"7f"),
  2150 => (x"08",x"1c",x"1c",x"3e"),
  2151 => (x"18",x"10",x"00",x"08"),
  2152 => (x"10",x"18",x"7c",x"7c"),
  2153 => (x"30",x"10",x"00",x"00"),
  2154 => (x"10",x"30",x"7c",x"7c"),
  2155 => (x"60",x"30",x"10",x"00"),
  2156 => (x"06",x"1e",x"78",x"60"),
  2157 => (x"3c",x"66",x"42",x"00"),
  2158 => (x"42",x"66",x"3c",x"18"),
  2159 => (x"6a",x"38",x"78",x"00"),
  2160 => (x"38",x"6c",x"c6",x"c2"),
  2161 => (x"00",x"00",x"60",x"00"),
  2162 => (x"60",x"00",x"00",x"60"),
  2163 => (x"5b",x"5e",x"0e",x"00"),
  2164 => (x"1e",x"0e",x"5d",x"5c"),
  2165 => (x"e7",x"c2",x"4c",x"71"),
  2166 => (x"c0",x"4d",x"bf",x"ce"),
  2167 => (x"74",x"1e",x"c0",x"4b"),
  2168 => (x"87",x"c7",x"02",x"ab"),
  2169 => (x"c0",x"48",x"a6",x"c4"),
  2170 => (x"c4",x"87",x"c5",x"78"),
  2171 => (x"78",x"c1",x"48",x"a6"),
  2172 => (x"73",x"1e",x"66",x"c4"),
  2173 => (x"87",x"db",x"ed",x"49"),
  2174 => (x"e0",x"c0",x"86",x"c8"),
  2175 => (x"87",x"cc",x"ef",x"49"),
  2176 => (x"6a",x"4a",x"a5",x"c4"),
  2177 => (x"87",x"ce",x"f0",x"49"),
  2178 => (x"cb",x"87",x"e4",x"f0"),
  2179 => (x"c8",x"83",x"c1",x"85"),
  2180 => (x"ff",x"04",x"ab",x"b7"),
  2181 => (x"26",x"26",x"87",x"c7"),
  2182 => (x"26",x"4c",x"26",x"4d"),
  2183 => (x"1e",x"4f",x"26",x"4b"),
  2184 => (x"e7",x"c2",x"4a",x"71"),
  2185 => (x"e7",x"c2",x"5a",x"d2"),
  2186 => (x"78",x"c7",x"48",x"d2"),
  2187 => (x"87",x"dd",x"fe",x"49"),
  2188 => (x"c1",x"1e",x"4f",x"26"),
  2189 => (x"ea",x"eb",x"49",x"c0"),
  2190 => (x"e2",x"d2",x"c2",x"87"),
  2191 => (x"26",x"78",x"c0",x"48"),
  2192 => (x"5b",x"5e",x"0e",x"4f"),
  2193 => (x"f4",x"0e",x"5d",x"5c"),
  2194 => (x"c8",x"7e",x"c0",x"86"),
  2195 => (x"bf",x"ec",x"48",x"a6"),
  2196 => (x"c2",x"80",x"fc",x"78"),
  2197 => (x"78",x"bf",x"ce",x"e7"),
  2198 => (x"bf",x"d6",x"e7",x"c2"),
  2199 => (x"4c",x"bf",x"e8",x"4d"),
  2200 => (x"c9",x"e7",x"49",x"c7"),
  2201 => (x"c2",x"49",x"70",x"87"),
  2202 => (x"87",x"d0",x"05",x"99"),
  2203 => (x"bf",x"da",x"d2",x"c2"),
  2204 => (x"c8",x"b9",x"ff",x"49"),
  2205 => (x"99",x"c1",x"99",x"66"),
  2206 => (x"87",x"eb",x"c0",x"02"),
  2207 => (x"ed",x"e6",x"49",x"c7"),
  2208 => (x"02",x"98",x"70",x"87"),
  2209 => (x"db",x"e2",x"87",x"cd"),
  2210 => (x"e6",x"49",x"c7",x"87"),
  2211 => (x"98",x"70",x"87",x"e0"),
  2212 => (x"c2",x"87",x"f3",x"05"),
  2213 => (x"4a",x"bf",x"e2",x"d2"),
  2214 => (x"d2",x"c2",x"ba",x"c1"),
  2215 => (x"c0",x"c1",x"5a",x"e6"),
  2216 => (x"fe",x"e9",x"49",x"a2"),
  2217 => (x"c2",x"7e",x"c1",x"87"),
  2218 => (x"c8",x"48",x"da",x"d2"),
  2219 => (x"d2",x"c2",x"78",x"66"),
  2220 => (x"c1",x"05",x"bf",x"e2"),
  2221 => (x"c0",x"c8",x"87",x"cb"),
  2222 => (x"d2",x"c2",x"7e",x"c0"),
  2223 => (x"49",x"13",x"4b",x"ca"),
  2224 => (x"70",x"87",x"eb",x"e5"),
  2225 => (x"87",x"c2",x"02",x"98"),
  2226 => (x"48",x"6e",x"b4",x"6e"),
  2227 => (x"c4",x"28",x"b7",x"c1"),
  2228 => (x"98",x"70",x"58",x"a6"),
  2229 => (x"87",x"e6",x"ff",x"05"),
  2230 => (x"ff",x"c3",x"49",x"74"),
  2231 => (x"c0",x"1e",x"71",x"99"),
  2232 => (x"87",x"f2",x"e7",x"49"),
  2233 => (x"b7",x"c8",x"49",x"74"),
  2234 => (x"c1",x"1e",x"71",x"29"),
  2235 => (x"87",x"e6",x"e7",x"49"),
  2236 => (x"fd",x"c3",x"86",x"c8"),
  2237 => (x"87",x"f6",x"e4",x"49"),
  2238 => (x"e4",x"49",x"fa",x"c3"),
  2239 => (x"c4",x"c6",x"87",x"f0"),
  2240 => (x"c3",x"49",x"74",x"87"),
  2241 => (x"b7",x"c8",x"99",x"ff"),
  2242 => (x"74",x"b4",x"71",x"2c"),
  2243 => (x"e2",x"c0",x"02",x"9c"),
  2244 => (x"48",x"a6",x"c8",x"87"),
  2245 => (x"78",x"bf",x"c8",x"ff"),
  2246 => (x"c2",x"49",x"66",x"c8"),
  2247 => (x"89",x"bf",x"de",x"d2"),
  2248 => (x"03",x"a9",x"c0",x"c2"),
  2249 => (x"4c",x"c0",x"87",x"c4"),
  2250 => (x"d2",x"c2",x"87",x"cf"),
  2251 => (x"66",x"c8",x"48",x"de"),
  2252 => (x"c2",x"87",x"c6",x"78"),
  2253 => (x"c0",x"48",x"de",x"d2"),
  2254 => (x"c8",x"49",x"74",x"78"),
  2255 => (x"87",x"ce",x"05",x"99"),
  2256 => (x"e3",x"49",x"f5",x"c3"),
  2257 => (x"49",x"70",x"87",x"e8"),
  2258 => (x"c0",x"02",x"99",x"c2"),
  2259 => (x"e7",x"c2",x"87",x"e6"),
  2260 => (x"c9",x"02",x"bf",x"d2"),
  2261 => (x"88",x"c1",x"48",x"87"),
  2262 => (x"58",x"d6",x"e7",x"c2"),
  2263 => (x"66",x"c4",x"87",x"d4"),
  2264 => (x"80",x"d8",x"c1",x"48"),
  2265 => (x"6e",x"58",x"a6",x"c4"),
  2266 => (x"c5",x"c0",x"02",x"bf"),
  2267 => (x"49",x"ff",x"4b",x"87"),
  2268 => (x"7e",x"c1",x"0f",x"73"),
  2269 => (x"99",x"c4",x"49",x"74"),
  2270 => (x"c3",x"87",x"ce",x"05"),
  2271 => (x"ed",x"e2",x"49",x"f2"),
  2272 => (x"c2",x"49",x"70",x"87"),
  2273 => (x"ee",x"c0",x"02",x"99"),
  2274 => (x"d2",x"e7",x"c2",x"87"),
  2275 => (x"48",x"6e",x"7e",x"bf"),
  2276 => (x"03",x"a8",x"b7",x"c7"),
  2277 => (x"6e",x"87",x"ca",x"c0"),
  2278 => (x"c2",x"80",x"c1",x"48"),
  2279 => (x"d4",x"58",x"d6",x"e7"),
  2280 => (x"48",x"66",x"c4",x"87"),
  2281 => (x"c4",x"80",x"d8",x"c1"),
  2282 => (x"bf",x"6e",x"58",x"a6"),
  2283 => (x"87",x"c5",x"c0",x"02"),
  2284 => (x"73",x"49",x"fe",x"4b"),
  2285 => (x"c3",x"7e",x"c1",x"0f"),
  2286 => (x"f1",x"e1",x"49",x"fd"),
  2287 => (x"c2",x"49",x"70",x"87"),
  2288 => (x"e3",x"c0",x"02",x"99"),
  2289 => (x"d2",x"e7",x"c2",x"87"),
  2290 => (x"c9",x"c0",x"02",x"bf"),
  2291 => (x"d2",x"e7",x"c2",x"87"),
  2292 => (x"c0",x"78",x"c0",x"48"),
  2293 => (x"66",x"c4",x"87",x"d0"),
  2294 => (x"82",x"d8",x"c1",x"4a"),
  2295 => (x"c5",x"c0",x"02",x"6a"),
  2296 => (x"49",x"fd",x"4b",x"87"),
  2297 => (x"7e",x"c1",x"0f",x"73"),
  2298 => (x"e1",x"49",x"fa",x"c3"),
  2299 => (x"49",x"70",x"87",x"c0"),
  2300 => (x"c0",x"02",x"99",x"c2"),
  2301 => (x"e7",x"c2",x"87",x"eb"),
  2302 => (x"c7",x"48",x"bf",x"d2"),
  2303 => (x"c0",x"03",x"a8",x"b7"),
  2304 => (x"e7",x"c2",x"87",x"c9"),
  2305 => (x"78",x"c7",x"48",x"d2"),
  2306 => (x"c4",x"87",x"d4",x"c0"),
  2307 => (x"d8",x"c1",x"48",x"66"),
  2308 => (x"58",x"a6",x"c4",x"80"),
  2309 => (x"c0",x"02",x"bf",x"6e"),
  2310 => (x"fc",x"4b",x"87",x"c5"),
  2311 => (x"c1",x"0f",x"73",x"49"),
  2312 => (x"c3",x"49",x"74",x"7e"),
  2313 => (x"c0",x"05",x"99",x"f0"),
  2314 => (x"da",x"c1",x"87",x"cf"),
  2315 => (x"fd",x"df",x"ff",x"49"),
  2316 => (x"c2",x"49",x"70",x"87"),
  2317 => (x"d0",x"c0",x"02",x"99"),
  2318 => (x"d2",x"e7",x"c2",x"87"),
  2319 => (x"cb",x"4b",x"49",x"bf"),
  2320 => (x"83",x"66",x"c4",x"93"),
  2321 => (x"73",x"71",x"4b",x"6b"),
  2322 => (x"02",x"9d",x"75",x"0f"),
  2323 => (x"6d",x"87",x"e9",x"c0"),
  2324 => (x"87",x"e4",x"c0",x"02"),
  2325 => (x"df",x"ff",x"49",x"6d"),
  2326 => (x"49",x"70",x"87",x"d4"),
  2327 => (x"c0",x"02",x"99",x"c1"),
  2328 => (x"a5",x"c4",x"87",x"cb"),
  2329 => (x"d2",x"e7",x"c2",x"4b"),
  2330 => (x"4b",x"6b",x"49",x"bf"),
  2331 => (x"02",x"85",x"c8",x"0f"),
  2332 => (x"6d",x"87",x"c5",x"c0"),
  2333 => (x"87",x"dc",x"ff",x"05"),
  2334 => (x"c8",x"c0",x"02",x"6e"),
  2335 => (x"d2",x"e7",x"c2",x"87"),
  2336 => (x"c8",x"f5",x"49",x"bf"),
  2337 => (x"f6",x"8e",x"f4",x"87"),
  2338 => (x"12",x"58",x"87",x"cd"),
  2339 => (x"1b",x"1d",x"14",x"11"),
  2340 => (x"59",x"5a",x"23",x"1c"),
  2341 => (x"f2",x"f5",x"94",x"91"),
  2342 => (x"00",x"00",x"f4",x"eb"),
  2343 => (x"00",x"00",x"00",x"00"),
  2344 => (x"00",x"00",x"00",x"00"),
  2345 => (x"19",x"a3",x"00",x"00"),
  2346 => (x"19",x"a3",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

