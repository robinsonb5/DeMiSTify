library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e4e8c287",
    12 => x"48c0c44e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90588",
    17 => x"49e4e8c2",
    18 => x"48f0d3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"f0d3c287",
    25 => x"ecd3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e0c187f7",
    29 => x"d3c287fc",
    30 => x"d3c24df0",
    31 => x"ad744cf0",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"c04b710e",
    37 => x"9a4a134c",
    38 => x"7287cd02",
    39 => x"87e0c049",
    40 => x"4a1384c1",
    41 => x"87f3059a",
    42 => x"4c264874",
    43 => x"4f264b26",
    44 => x"8148731e",
    45 => x"c502a973",
    46 => x"05531287",
    47 => x"4f2687f6",
    48 => x"c0ff1e1e",
    49 => x"c4486a4a",
    50 => x"a6c498c0",
    51 => x"02987058",
    52 => x"7a7187f3",
    53 => x"4f262648",
    54 => x"ff1e731e",
    55 => x"ffc34bd4",
    56 => x"c34a6b7b",
    57 => x"496b7bff",
    58 => x"b17232c8",
    59 => x"6b7bffc3",
    60 => x"7131c84a",
    61 => x"7bffc3b2",
    62 => x"32c8496b",
    63 => x"4871b172",
    64 => x"4d2687c4",
    65 => x"4b264c26",
    66 => x"5e0e4f26",
    67 => x"0e5d5c5b",
    68 => x"d4ff4a71",
    69 => x"c348724c",
    70 => x"7c7098ff",
    71 => x"bff0d3c2",
    72 => x"d087c805",
    73 => x"30c94866",
    74 => x"d058a6d4",
    75 => x"29d84966",
    76 => x"ffc34871",
    77 => x"d07c7098",
    78 => x"29d04966",
    79 => x"ffc34871",
    80 => x"d07c7098",
    81 => x"29c84966",
    82 => x"ffc34871",
    83 => x"d07c7098",
    84 => x"ffc34866",
    85 => x"727c7098",
    86 => x"7129d049",
    87 => x"98ffc348",
    88 => x"4b6c7c70",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87fffd",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487dffd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c1fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87defc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"49e3c878",
   125 => x"d387d5fa",
   126 => x"c01ec04b",
   127 => x"c1c1f0ff",
   128 => x"87c6fc49",
   129 => x"987086c4",
   130 => x"ff87ca05",
   131 => x"ffc348d4",
   132 => x"cb48c178",
   133 => x"87ebfd87",
   134 => x"ff058bc1",
   135 => x"48c087db",
   136 => x"4387e3fb",
   137 => x"5300444d",
   138 => x"20434844",
   139 => x"6c696166",
   140 => x"49000a21",
   141 => x"00525245",
   142 => x"00495053",
   143 => x"74697257",
   144 => x"61662065",
   145 => x"64656c69",
   146 => x"5e0e000a",
   147 => x"ff0e5c5b",
   148 => x"eefc4cd4",
   149 => x"1eeac687",
   150 => x"c1f0e1c0",
   151 => x"e9fa49c8",
   152 => x"c186c487",
   153 => x"87c802a8",
   154 => x"c087fdfd",
   155 => x"87e8c148",
   156 => x"7087e5f9",
   157 => x"ffffcf49",
   158 => x"a9eac699",
   159 => x"fd87c802",
   160 => x"48c087e6",
   161 => x"c387d1c1",
   162 => x"f1c07cff",
   163 => x"87c7fc4b",
   164 => x"c0029870",
   165 => x"1ec087eb",
   166 => x"c1f0ffc0",
   167 => x"e9f949fa",
   168 => x"7086c487",
   169 => x"87d90598",
   170 => x"6c7cffc3",
   171 => x"7cffc349",
   172 => x"c17c7c7c",
   173 => x"c40299c0",
   174 => x"db48c187",
   175 => x"d748c087",
   176 => x"05abc287",
   177 => x"e7c887ca",
   178 => x"87c0f749",
   179 => x"87c848c0",
   180 => x"fe058bc1",
   181 => x"48c087f7",
   182 => x"0e87e9f8",
   183 => x"5d5c5b5e",
   184 => x"d0ff1e0e",
   185 => x"c0c0c84d",
   186 => x"f0d3c24b",
   187 => x"c878c148",
   188 => x"d7f649f8",
   189 => x"6d4cc787",
   190 => x"c4987348",
   191 => x"987058a6",
   192 => x"6d87cc02",
   193 => x"c4987348",
   194 => x"987058a6",
   195 => x"c287f405",
   196 => x"87eff97d",
   197 => x"9873486d",
   198 => x"7058a6c4",
   199 => x"87cc0298",
   200 => x"9873486d",
   201 => x"7058a6c4",
   202 => x"87f40598",
   203 => x"1ec07dc3",
   204 => x"c1d0e5c0",
   205 => x"d1f749c0",
   206 => x"c186c487",
   207 => x"87c105a8",
   208 => x"05acc24c",
   209 => x"f3c887cb",
   210 => x"87c0f549",
   211 => x"cec148c0",
   212 => x"058cc187",
   213 => x"fb87e0fe",
   214 => x"d3c287f0",
   215 => x"987058f4",
   216 => x"c187cd05",
   217 => x"f0ffc01e",
   218 => x"f649d0c1",
   219 => x"86c487dc",
   220 => x"c348d4ff",
   221 => x"ddc578ff",
   222 => x"f8d3c287",
   223 => x"73486d58",
   224 => x"58a6c498",
   225 => x"cc029870",
   226 => x"73486d87",
   227 => x"58a6c498",
   228 => x"f4059870",
   229 => x"ff7dc287",
   230 => x"ffc348d4",
   231 => x"2648c178",
   232 => x"0e87dff5",
   233 => x"5d5c5b5e",
   234 => x"c0c81e0e",
   235 => x"4cc04bc0",
   236 => x"dfcdeec5",
   237 => x"5ca6c44a",
   238 => x"c34cd4ff",
   239 => x"486c7cff",
   240 => x"05a8fec3",
   241 => x"7187c0c2",
   242 => x"e2c00599",
   243 => x"bfd0ff87",
   244 => x"c4987348",
   245 => x"987058a6",
   246 => x"ff87ce02",
   247 => x"7348bfd0",
   248 => x"58a6c498",
   249 => x"f2059870",
   250 => x"48d0ff87",
   251 => x"d478d1c4",
   252 => x"b7c04866",
   253 => x"e0c006a8",
   254 => x"7cffc387",
   255 => x"99714a6c",
   256 => x"7187c702",
   257 => x"0a7a970a",
   258 => x"66d481c1",
   259 => x"d888c148",
   260 => x"b7c058a6",
   261 => x"e0ff01a8",
   262 => x"7cffc387",
   263 => x"0599717c",
   264 => x"ff87e1c0",
   265 => x"7348bfd0",
   266 => x"58a6c498",
   267 => x"ce029870",
   268 => x"bfd0ff87",
   269 => x"c4987348",
   270 => x"987058a6",
   271 => x"ff87f205",
   272 => x"78d048d0",
   273 => x"c17e4ac1",
   274 => x"eefd058a",
   275 => x"26486e87",
   276 => x"0e87eff2",
   277 => x"0e5c5b5e",
   278 => x"c84a711e",
   279 => x"c04bc0c0",
   280 => x"48d4ff4c",
   281 => x"ff78ffc3",
   282 => x"7348bfd0",
   283 => x"58a6c498",
   284 => x"ce029870",
   285 => x"bfd0ff87",
   286 => x"c4987348",
   287 => x"987058a6",
   288 => x"ff87f205",
   289 => x"c3c448d0",
   290 => x"48d4ff78",
   291 => x"7278ffc3",
   292 => x"f0ffc01e",
   293 => x"f149d1c1",
   294 => x"86c487f0",
   295 => x"c0059870",
   296 => x"c0c887ee",
   297 => x"4966d41e",
   298 => x"c487f8fb",
   299 => x"ff4c7086",
   300 => x"7348bfd0",
   301 => x"58a6c498",
   302 => x"ce029870",
   303 => x"bfd0ff87",
   304 => x"c4987348",
   305 => x"987058a6",
   306 => x"ff87f205",
   307 => x"78c248d0",
   308 => x"f0264874",
   309 => x"5e0e87ee",
   310 => x"0e5d5c5b",
   311 => x"ffc01ec0",
   312 => x"49c9c1f0",
   313 => x"d287e3f0",
   314 => x"fed3c21e",
   315 => x"87f3fa49",
   316 => x"4cc086c8",
   317 => x"b7d284c1",
   318 => x"87f804ac",
   319 => x"97fed3c2",
   320 => x"c0c349bf",
   321 => x"a9c0c199",
   322 => x"87e7c005",
   323 => x"97c5d4c2",
   324 => x"31d049bf",
   325 => x"97c6d4c2",
   326 => x"32c84abf",
   327 => x"d4c2b172",
   328 => x"4abf97c7",
   329 => x"cf4c71b1",
   330 => x"9cffffff",
   331 => x"34ca84c1",
   332 => x"c287e7c1",
   333 => x"bf97c7d4",
   334 => x"c631c149",
   335 => x"c8d4c299",
   336 => x"c74abf97",
   337 => x"b1722ab7",
   338 => x"97c3d4c2",
   339 => x"cf4d4abf",
   340 => x"c4d4c29d",
   341 => x"c34abf97",
   342 => x"c232ca9a",
   343 => x"bf97c5d4",
   344 => x"7333c24b",
   345 => x"c6d4c2b2",
   346 => x"c34bbf97",
   347 => x"b7c69bc0",
   348 => x"c2b2732b",
   349 => x"7148c181",
   350 => x"c1497030",
   351 => x"70307548",
   352 => x"c14c724d",
   353 => x"c8947184",
   354 => x"06adb7c0",
   355 => x"34c187cc",
   356 => x"c0c82db7",
   357 => x"ff01adb7",
   358 => x"487487f4",
   359 => x"0e87e3ed",
   360 => x"0e5c5b5e",
   361 => x"4cc04b71",
   362 => x"c04866d0",
   363 => x"c006a8b7",
   364 => x"4a1387e3",
   365 => x"bf9766cc",
   366 => x"4866cc49",
   367 => x"a6d080c1",
   368 => x"aab77158",
   369 => x"c187c402",
   370 => x"c187cc48",
   371 => x"b766d084",
   372 => x"ddff04ac",
   373 => x"c248c087",
   374 => x"264d2687",
   375 => x"264b264c",
   376 => x"5b5e0e4f",
   377 => x"c20e5d5c",
   378 => x"c048e4dc",
   379 => x"dcd4c278",
   380 => x"f949c01e",
   381 => x"86c487dd",
   382 => x"c5059870",
   383 => x"c848c087",
   384 => x"4bc087ef",
   385 => x"48dce1c2",
   386 => x"1ec878c1",
   387 => x"1efde0c0",
   388 => x"49d2d5c2",
   389 => x"c887c8fe",
   390 => x"05987086",
   391 => x"e1c287c6",
   392 => x"78c048dc",
   393 => x"e1c01ec8",
   394 => x"d5c21ec6",
   395 => x"eefd49ee",
   396 => x"7086c887",
   397 => x"87c60598",
   398 => x"48dce1c2",
   399 => x"e1c278c0",
   400 => x"c002bfdc",
   401 => x"dbc287fa",
   402 => x"c24bbfe2",
   403 => x"bf9fdadc",
   404 => x"ead6c54a",
   405 => x"87c705aa",
   406 => x"bfe2dbc2",
   407 => x"ca87cc4b",
   408 => x"02aad5e9",
   409 => x"48c087c5",
   410 => x"c287c6c7",
   411 => x"731edcd4",
   412 => x"87dff749",
   413 => x"987086c4",
   414 => x"c087c505",
   415 => x"87f1c648",
   416 => x"e1c01ec8",
   417 => x"d5c21ecf",
   418 => x"d2fc49ee",
   419 => x"7086c887",
   420 => x"87c80598",
   421 => x"48e4dcc2",
   422 => x"87da78c1",
   423 => x"e1c01ec8",
   424 => x"d5c21ed8",
   425 => x"f6fb49d2",
   426 => x"7086c887",
   427 => x"c5c00298",
   428 => x"c548c087",
   429 => x"dcc287fb",
   430 => x"49bf97da",
   431 => x"05a9d5c1",
   432 => x"c287cdc0",
   433 => x"bf97dbdc",
   434 => x"a9eac249",
   435 => x"87c5c002",
   436 => x"dcc548c0",
   437 => x"dcd4c287",
   438 => x"c34cbf97",
   439 => x"c002ace9",
   440 => x"ebc387cc",
   441 => x"c5c002ac",
   442 => x"c548c087",
   443 => x"d4c287c3",
   444 => x"49bf97e7",
   445 => x"ccc00599",
   446 => x"e8d4c287",
   447 => x"c249bf97",
   448 => x"c5c002a9",
   449 => x"c448c087",
   450 => x"d4c287e7",
   451 => x"48bf97e9",
   452 => x"58e0dcc2",
   453 => x"dcc288c1",
   454 => x"d4c258e4",
   455 => x"49bf97ea",
   456 => x"d4c28173",
   457 => x"4abf97eb",
   458 => x"7135c84d",
   459 => x"fce0c285",
   460 => x"ecd4c25d",
   461 => x"c248bf97",
   462 => x"c258d0e1",
   463 => x"02bfe4dc",
   464 => x"c887dcc2",
   465 => x"f4e0c01e",
   466 => x"eed5c21e",
   467 => x"87cff949",
   468 => x"987086c8",
   469 => x"87c5c002",
   470 => x"d4c348c0",
   471 => x"dcdcc287",
   472 => x"c4484abf",
   473 => x"ecdcc230",
   474 => x"cce1c258",
   475 => x"c1d5c25a",
   476 => x"c849bf97",
   477 => x"c0d5c231",
   478 => x"a14bbf97",
   479 => x"c2d5c249",
   480 => x"d04bbf97",
   481 => x"49a17333",
   482 => x"97c3d5c2",
   483 => x"33d84bbf",
   484 => x"c249a173",
   485 => x"c259d4e1",
   486 => x"91bfcce1",
   487 => x"bff8e0c2",
   488 => x"c0e1c281",
   489 => x"c9d5c259",
   490 => x"c84bbf97",
   491 => x"c8d5c233",
   492 => x"a34cbf97",
   493 => x"cad5c24b",
   494 => x"d04cbf97",
   495 => x"4ba37434",
   496 => x"97cbd5c2",
   497 => x"9ccf4cbf",
   498 => x"a37434d8",
   499 => x"c4e1c24b",
   500 => x"738bc25b",
   501 => x"c4e1c292",
   502 => x"78a17248",
   503 => x"c287cbc1",
   504 => x"bf97eed4",
   505 => x"c231c849",
   506 => x"bf97edd4",
   507 => x"c249a14a",
   508 => x"c559ecdc",
   509 => x"81ffc731",
   510 => x"e1c229c9",
   511 => x"d4c259cc",
   512 => x"4abf97f3",
   513 => x"d4c232c8",
   514 => x"4bbf97f2",
   515 => x"e1c24aa2",
   516 => x"e1c25ad4",
   517 => x"7592bfcc",
   518 => x"c8e1c282",
   519 => x"c0e1c25a",
   520 => x"c278c048",
   521 => x"7248fce0",
   522 => x"49c078a1",
   523 => x"c187f7c7",
   524 => x"87e5f648",
   525 => x"33544146",
   526 => x"20202032",
   527 => x"54414600",
   528 => x"20203631",
   529 => x"41460020",
   530 => x"20323354",
   531 => x"46002020",
   532 => x"32335441",
   533 => x"00202020",
   534 => x"31544146",
   535 => x"20202036",
   536 => x"5b5e0e00",
   537 => x"710e5d5c",
   538 => x"e4dcc24a",
   539 => x"87cc02bf",
   540 => x"b7c74b72",
   541 => x"c14d722b",
   542 => x"87ca9dff",
   543 => x"b7c84b72",
   544 => x"c34d722b",
   545 => x"d4c29dff",
   546 => x"e0c21edc",
   547 => x"7349bff8",
   548 => x"feee7181",
   549 => x"7086c487",
   550 => x"87c50598",
   551 => x"e6c048c0",
   552 => x"e4dcc287",
   553 => x"87d202bf",
   554 => x"91c44975",
   555 => x"81dcd4c2",
   556 => x"ffcf4c69",
   557 => x"9cffffff",
   558 => x"497587cb",
   559 => x"d4c291c2",
   560 => x"699f81dc",
   561 => x"f448744c",
   562 => x"5e0e87cf",
   563 => x"0e5d5c5b",
   564 => x"4c7186f4",
   565 => x"e1c24bc0",
   566 => x"c47ebfd4",
   567 => x"e1c248a6",
   568 => x"c878bfd8",
   569 => x"78c048a6",
   570 => x"bfe8dcc2",
   571 => x"06a8c048",
   572 => x"c887ddc2",
   573 => x"99cf4966",
   574 => x"c287d805",
   575 => x"c81edcd4",
   576 => x"c1484966",
   577 => x"58a6cc80",
   578 => x"c487c8ed",
   579 => x"dcd4c286",
   580 => x"c087c34b",
   581 => x"6b9783e0",
   582 => x"c1029a4a",
   583 => x"e5c387e1",
   584 => x"dac102aa",
   585 => x"49a3cb87",
   586 => x"d8496997",
   587 => x"cec10599",
   588 => x"c01ecb87",
   589 => x"731e66e0",
   590 => x"87e3f149",
   591 => x"987086c8",
   592 => x"87fbc005",
   593 => x"c44aa3dc",
   594 => x"796a49a4",
   595 => x"c849a3da",
   596 => x"699f4da4",
   597 => x"dcc27d48",
   598 => x"d302bfe4",
   599 => x"49a3d487",
   600 => x"c049699f",
   601 => x"7199ffff",
   602 => x"c430d048",
   603 => x"87c258a6",
   604 => x"486e7ec0",
   605 => x"7d70806d",
   606 => x"48c17cc0",
   607 => x"c887c5c1",
   608 => x"80c14866",
   609 => x"c258a6cc",
   610 => x"a8bfe8dc",
   611 => x"87e3fd04",
   612 => x"bfe4dcc2",
   613 => x"87eac002",
   614 => x"c4fb496e",
   615 => x"58a6c487",
   616 => x"ffcf4970",
   617 => x"99f8ffff",
   618 => x"87d602a9",
   619 => x"89c24970",
   620 => x"bfdcdcc2",
   621 => x"fce0c291",
   622 => x"807148bf",
   623 => x"fc58a6c8",
   624 => x"48c087e1",
   625 => x"d0f08ef4",
   626 => x"1e731e87",
   627 => x"496a4a71",
   628 => x"7a7181c1",
   629 => x"bfe0dcc2",
   630 => x"87cb0599",
   631 => x"6b4ba2c8",
   632 => x"87fdf949",
   633 => x"c17b4970",
   634 => x"87f1ef48",
   635 => x"711e731e",
   636 => x"fce0c24b",
   637 => x"a3c849bf",
   638 => x"c24a6a4a",
   639 => x"dcdcc28a",
   640 => x"a17292bf",
   641 => x"e0dcc249",
   642 => x"9a6b4abf",
   643 => x"c849a172",
   644 => x"e8711e66",
   645 => x"86c487fd",
   646 => x"c4059870",
   647 => x"c248c087",
   648 => x"ee48c187",
   649 => x"5e0e87f7",
   650 => x"710e5c5b",
   651 => x"724bc04a",
   652 => x"e0c0029a",
   653 => x"49a2da87",
   654 => x"c24b699f",
   655 => x"02bfe4dc",
   656 => x"a2d487cf",
   657 => x"49699f49",
   658 => x"ffffc04c",
   659 => x"c234d09c",
   660 => x"744cc087",
   661 => x"029b73b3",
   662 => x"c24a87df",
   663 => x"dcdcc28a",
   664 => x"c29249bf",
   665 => x"48bffce0",
   666 => x"e1c28072",
   667 => x"487158dc",
   668 => x"dcc230c4",
   669 => x"e9c058ec",
   670 => x"c0e1c287",
   671 => x"e1c24bbf",
   672 => x"e1c248d8",
   673 => x"c278bfc4",
   674 => x"02bfe4dc",
   675 => x"dcc287c9",
   676 => x"c449bfdc",
   677 => x"c287c731",
   678 => x"49bfc8e1",
   679 => x"dcc231c4",
   680 => x"e1c259ec",
   681 => x"f2ec5bd8",
   682 => x"5b5e0e87",
   683 => x"f40e5d5c",
   684 => x"9a4a7186",
   685 => x"c287de02",
   686 => x"c048d8d4",
   687 => x"d0d4c278",
   688 => x"d8e1c248",
   689 => x"d4c278bf",
   690 => x"e1c248d4",
   691 => x"c078bfd4",
   692 => x"c048fff1",
   693 => x"e8dcc278",
   694 => x"d4c249bf",
   695 => x"714abfd8",
   696 => x"cbc403aa",
   697 => x"cf497287",
   698 => x"e0c00599",
   699 => x"dcd4c287",
   700 => x"d0d4c21e",
   701 => x"d4c249bf",
   702 => x"a1c148d0",
   703 => x"d2e57178",
   704 => x"c086c487",
   705 => x"c248fbf1",
   706 => x"cc78dcd4",
   707 => x"fbf1c087",
   708 => x"e0c048bf",
   709 => x"fff1c080",
   710 => x"d8d4c258",
   711 => x"80c148bf",
   712 => x"58dcd4c2",
   713 => x"000c7b27",
   714 => x"bf97bf00",
   715 => x"c2029c4c",
   716 => x"e5c387ee",
   717 => x"e7c202ac",
   718 => x"fbf1c087",
   719 => x"a3cb4bbf",
   720 => x"cf4d1149",
   721 => x"d6c105ad",
   722 => x"df497487",
   723 => x"cd89c199",
   724 => x"ecdcc291",
   725 => x"4aa3c181",
   726 => x"a3c35112",
   727 => x"c551124a",
   728 => x"51124aa3",
   729 => x"124aa3c7",
   730 => x"4aa3c951",
   731 => x"a3ce5112",
   732 => x"d051124a",
   733 => x"51124aa3",
   734 => x"124aa3d2",
   735 => x"4aa3d451",
   736 => x"a3d65112",
   737 => x"d851124a",
   738 => x"51124aa3",
   739 => x"124aa3dc",
   740 => x"4aa3de51",
   741 => x"f1c05112",
   742 => x"78c148ff",
   743 => x"7587c1c1",
   744 => x"0599c849",
   745 => x"7587f3c0",
   746 => x"0599d049",
   747 => x"66dc87d0",
   748 => x"87cac002",
   749 => x"66dc4973",
   750 => x"0298700f",
   751 => x"f1c087dc",
   752 => x"c005bfff",
   753 => x"dcc287c6",
   754 => x"50c048ec",
   755 => x"48fff1c0",
   756 => x"f1c078c0",
   757 => x"c248bffb",
   758 => x"f1c087dc",
   759 => x"78c048ff",
   760 => x"bfe8dcc2",
   761 => x"d8d4c249",
   762 => x"aa714abf",
   763 => x"87f5fb04",
   764 => x"bfd8e1c2",
   765 => x"87c8c005",
   766 => x"bfe4dcc2",
   767 => x"87f4c102",
   768 => x"bfd4d4c2",
   769 => x"87d9f149",
   770 => x"58d8d4c2",
   771 => x"dcc27e70",
   772 => x"c002bfe4",
   773 => x"496e87dd",
   774 => x"ffffffcf",
   775 => x"02a999f8",
   776 => x"c487c8c0",
   777 => x"78c048a6",
   778 => x"c487e6c0",
   779 => x"78c148a6",
   780 => x"6e87dec0",
   781 => x"f8ffcf49",
   782 => x"c002a999",
   783 => x"a6c887c8",
   784 => x"c078c048",
   785 => x"a6c887c5",
   786 => x"c478c148",
   787 => x"66c848a6",
   788 => x"0566c478",
   789 => x"6e87ddc0",
   790 => x"c289c249",
   791 => x"91bfdcdc",
   792 => x"bffce0c2",
   793 => x"c2807148",
   794 => x"c258d4d4",
   795 => x"c048d8d4",
   796 => x"87e1f978",
   797 => x"8ef448c0",
   798 => x"0087dee5",
   799 => x"00000000",
   800 => x"1e000000",
   801 => x"c348d4ff",
   802 => x"496878ff",
   803 => x"87c60299",
   804 => x"05a9fbc0",
   805 => x"487187ee",
   806 => x"5e0e4f26",
   807 => x"710e5c5b",
   808 => x"ff4bc04a",
   809 => x"ffc348d4",
   810 => x"99496878",
   811 => x"87c1c102",
   812 => x"02a9ecc0",
   813 => x"c087fac0",
   814 => x"c002a9fb",
   815 => x"66cc87f3",
   816 => x"cc03abb7",
   817 => x"0266d087",
   818 => x"097287c7",
   819 => x"c1097997",
   820 => x"02997182",
   821 => x"83c187c2",
   822 => x"c348d4ff",
   823 => x"496878ff",
   824 => x"87cd0299",
   825 => x"02a9ecc0",
   826 => x"fbc087c7",
   827 => x"cdff05a9",
   828 => x"0266d087",
   829 => x"97c087c3",
   830 => x"a9fbc07a",
   831 => x"7387c705",
   832 => x"8c0cc04c",
   833 => x"4c7387c2",
   834 => x"87c24874",
   835 => x"4c264d26",
   836 => x"4f264b26",
   837 => x"48d4ff1e",
   838 => x"6878ffc3",
   839 => x"b7f0c049",
   840 => x"87ca04a9",
   841 => x"a9b7f9c0",
   842 => x"c087c301",
   843 => x"c1c189f0",
   844 => x"ca04a9b7",
   845 => x"b7c6c187",
   846 => x"87c301a9",
   847 => x"7189f7c0",
   848 => x"0e4f2648",
   849 => x"5d5c5b5e",
   850 => x"7186f40e",
   851 => x"4bd4ff4c",
   852 => x"c37e4dc0",
   853 => x"d0ff7bff",
   854 => x"c0c848bf",
   855 => x"a6c898c0",
   856 => x"02987058",
   857 => x"d0ff87d0",
   858 => x"c0c848bf",
   859 => x"a6c898c0",
   860 => x"05987058",
   861 => x"d0ff87f0",
   862 => x"78e1c048",
   863 => x"c2fc7bd4",
   864 => x"99497087",
   865 => x"87c7c102",
   866 => x"c87bffc3",
   867 => x"786b48a6",
   868 => x"c04866c8",
   869 => x"c802a8fb",
   870 => x"f4e1c287",
   871 => x"eec002bf",
   872 => x"714dc187",
   873 => x"e6c00299",
   874 => x"a9fbc087",
   875 => x"fb87c302",
   876 => x"ffc387d1",
   877 => x"c1496b7b",
   878 => x"cc05a9c6",
   879 => x"7bffc387",
   880 => x"48a6c87b",
   881 => x"49c0786b",
   882 => x"0599714d",
   883 => x"7587daff",
   884 => x"dec1059d",
   885 => x"7bffc387",
   886 => x"ffc34a6b",
   887 => x"48a6c47b",
   888 => x"486e786b",
   889 => x"a6c480c1",
   890 => x"49a4c858",
   891 => x"c8496997",
   892 => x"da05a966",
   893 => x"49a4c987",
   894 => x"aa496997",
   895 => x"ca87d005",
   896 => x"699749a4",
   897 => x"a966c449",
   898 => x"c187c405",
   899 => x"c887d64d",
   900 => x"ecc04866",
   901 => x"87c902a8",
   902 => x"c04866c8",
   903 => x"c405a8fb",
   904 => x"c17ec087",
   905 => x"7bffc34d",
   906 => x"6b48a6c8",
   907 => x"029d7578",
   908 => x"ff87e2fe",
   909 => x"c848bfd0",
   910 => x"c898c0c0",
   911 => x"987058a6",
   912 => x"ff87d002",
   913 => x"c848bfd0",
   914 => x"c898c0c0",
   915 => x"987058a6",
   916 => x"ff87f005",
   917 => x"e0c048d0",
   918 => x"f4486e78",
   919 => x"87ecfa8e",
   920 => x"5c5b5e0e",
   921 => x"86f40e5d",
   922 => x"ff59a6c4",
   923 => x"c0c84cd0",
   924 => x"1e6e4bc0",
   925 => x"49f8e1c2",
   926 => x"c487cfe9",
   927 => x"02987086",
   928 => x"c287f7c5",
   929 => x"4dbffce1",
   930 => x"f6fa496e",
   931 => x"58a6c887",
   932 => x"9873486c",
   933 => x"7058a6cc",
   934 => x"87cc0298",
   935 => x"9873486c",
   936 => x"7058a6c4",
   937 => x"87f40598",
   938 => x"d4ff7cc5",
   939 => x"78d5c148",
   940 => x"bff4e1c2",
   941 => x"c481c149",
   942 => x"8ac14a66",
   943 => x"487232c6",
   944 => x"d4ffb071",
   945 => x"486c7808",
   946 => x"a6c49873",
   947 => x"02987058",
   948 => x"486c87cc",
   949 => x"a6c49873",
   950 => x"05987058",
   951 => x"7cc487f4",
   952 => x"c348d4ff",
   953 => x"486c78ff",
   954 => x"a6c49873",
   955 => x"02987058",
   956 => x"486c87cc",
   957 => x"a6c49873",
   958 => x"05987058",
   959 => x"7cc587f4",
   960 => x"c148d4ff",
   961 => x"78c178d3",
   962 => x"9873486c",
   963 => x"7058a6c4",
   964 => x"87cc0298",
   965 => x"9873486c",
   966 => x"7058a6c4",
   967 => x"87f40598",
   968 => x"9d757cc4",
   969 => x"87d0c202",
   970 => x"7edcd4c2",
   971 => x"f8e1c21e",
   972 => x"87f8ea49",
   973 => x"987086c4",
   974 => x"c087c505",
   975 => x"87fcc248",
   976 => x"adb7c0c8",
   977 => x"4a87c404",
   978 => x"7587c48d",
   979 => x"6c4dc04a",
   980 => x"c8987348",
   981 => x"987058a6",
   982 => x"6c87cc02",
   983 => x"c8987348",
   984 => x"987058a6",
   985 => x"cd87f405",
   986 => x"48d4ff7c",
   987 => x"7278d4c1",
   988 => x"718ac149",
   989 => x"87d90299",
   990 => x"48bf976e",
   991 => x"7808d4ff",
   992 => x"80c1486e",
   993 => x"7258a6c4",
   994 => x"718ac149",
   995 => x"e7ff0599",
   996 => x"73486c87",
   997 => x"58a6c498",
   998 => x"cc029870",
   999 => x"73486c87",
  1000 => x"58a6c498",
  1001 => x"f4059870",
  1002 => x"c27cc487",
  1003 => x"e849f8e1",
  1004 => x"9d7587d7",
  1005 => x"87f0fd05",
  1006 => x"9873486c",
  1007 => x"7058a6c4",
  1008 => x"87cd0298",
  1009 => x"9873486c",
  1010 => x"7058a6c4",
  1011 => x"f3ff0598",
  1012 => x"ff7cc587",
  1013 => x"d3c148d4",
  1014 => x"6c78c078",
  1015 => x"c4987348",
  1016 => x"987058a6",
  1017 => x"6c87cd02",
  1018 => x"c4987348",
  1019 => x"987058a6",
  1020 => x"87f3ff05",
  1021 => x"48c17cc4",
  1022 => x"48c087c2",
  1023 => x"cbf48ef4",
  1024 => x"5b5e0e87",
  1025 => x"1e0e5d5c",
  1026 => x"4cc04b71",
  1027 => x"04abb74d",
  1028 => x"c087e9c0",
  1029 => x"751ec3f5",
  1030 => x"87c4029d",
  1031 => x"87c24ac0",
  1032 => x"49724ac1",
  1033 => x"c487c2ea",
  1034 => x"c158a686",
  1035 => x"c2056e84",
  1036 => x"c14c7387",
  1037 => x"acb77385",
  1038 => x"87d7ff06",
  1039 => x"f326486e",
  1040 => x"5e0e87ca",
  1041 => x"0e5d5c5b",
  1042 => x"c2494c71",
  1043 => x"81bfcce2",
  1044 => x"7087eefe",
  1045 => x"c0029d4d",
  1046 => x"dcc287f3",
  1047 => x"4a754bec",
  1048 => x"c1ff49cb",
  1049 => x"4b7487ca",
  1050 => x"e4c193cb",
  1051 => x"83c483db",
  1052 => x"7bdac2c1",
  1053 => x"c5c14974",
  1054 => x"497487f6",
  1055 => x"e2c291de",
  1056 => x"807148e0",
  1057 => x"dcc27b70",
  1058 => x"d3f749ec",
  1059 => x"c1497487",
  1060 => x"c187ddc5",
  1061 => x"f187fec6",
  1062 => x"6f4c87f2",
  1063 => x"6e696461",
  1064 => x"2e2e2e67",
  1065 => x"42208000",
  1066 => x"006b6361",
  1067 => x"64616f4c",
  1068 => x"202e2a20",
  1069 => x"00203a00",
  1070 => x"61422080",
  1071 => x"80006b63",
  1072 => x"69784520",
  1073 => x"44530074",
  1074 => x"696e4920",
  1075 => x"002e2e74",
  1076 => x"42004b4f",
  1077 => x"20544f4f",
  1078 => x"52202020",
  1079 => x"1e004d4f",
  1080 => x"4b711e73",
  1081 => x"cce2c249",
  1082 => x"d4fc81bf",
  1083 => x"9a4a7087",
  1084 => x"4987c402",
  1085 => x"c287efe4",
  1086 => x"c048cce2",
  1087 => x"c1497378",
  1088 => x"cbf087f8",
  1089 => x"1e731e87",
  1090 => x"a3c44b71",
  1091 => x"d0c1024a",
  1092 => x"028ac187",
  1093 => x"028a87dc",
  1094 => x"8a87f2c0",
  1095 => x"87d3c105",
  1096 => x"bfcce2c2",
  1097 => x"87cbc102",
  1098 => x"c288c148",
  1099 => x"c158d0e2",
  1100 => x"e2c287c1",
  1101 => x"c649bfcc",
  1102 => x"d0e2c289",
  1103 => x"a9b7c059",
  1104 => x"87efc003",
  1105 => x"48cce2c2",
  1106 => x"e6c078c0",
  1107 => x"c8e2c287",
  1108 => x"87df02bf",
  1109 => x"bfcce2c2",
  1110 => x"c280c148",
  1111 => x"d258d0e2",
  1112 => x"c8e2c287",
  1113 => x"87cb02bf",
  1114 => x"bfcce2c2",
  1115 => x"c280c648",
  1116 => x"7358d0e2",
  1117 => x"ee87c349",
  1118 => x"5e0e87d6",
  1119 => x"0e5d5c5b",
  1120 => x"a6d086f0",
  1121 => x"dcd4c259",
  1122 => x"c24cc04d",
  1123 => x"c148c8e2",
  1124 => x"48a6c478",
  1125 => x"e2c278c0",
  1126 => x"c048bfcc",
  1127 => x"c106a8b7",
  1128 => x"d4c287c1",
  1129 => x"029848dc",
  1130 => x"c087f8c0",
  1131 => x"c81ec3f5",
  1132 => x"87c70266",
  1133 => x"c048a6c4",
  1134 => x"c487c578",
  1135 => x"78c148a6",
  1136 => x"e34966c4",
  1137 => x"86c487e3",
  1138 => x"84c14d70",
  1139 => x"c14866c4",
  1140 => x"58a6c880",
  1141 => x"bfcce2c2",
  1142 => x"c603acb7",
  1143 => x"059d7587",
  1144 => x"c087c8ff",
  1145 => x"029d754c",
  1146 => x"c087dec3",
  1147 => x"c81ec3f5",
  1148 => x"87c70266",
  1149 => x"c048a6cc",
  1150 => x"cc87c578",
  1151 => x"78c148a6",
  1152 => x"e24966cc",
  1153 => x"86c487e3",
  1154 => x"026e58a6",
  1155 => x"4987e6c2",
  1156 => x"699781cb",
  1157 => x"0299d049",
  1158 => x"c187d6c1",
  1159 => x"744adfc3",
  1160 => x"c191cb49",
  1161 => x"7281dbe4",
  1162 => x"c381c879",
  1163 => x"497451ff",
  1164 => x"e2c291de",
  1165 => x"85714de0",
  1166 => x"7d97c1c2",
  1167 => x"c049a5c1",
  1168 => x"dcc251e0",
  1169 => x"02bf97ec",
  1170 => x"84c187d2",
  1171 => x"c24ba5c2",
  1172 => x"db4aecdc",
  1173 => x"d7f9fe49",
  1174 => x"87d9c187",
  1175 => x"c049a5cd",
  1176 => x"c284c151",
  1177 => x"4a6e4ba5",
  1178 => x"f9fe49cb",
  1179 => x"c4c187c2",
  1180 => x"cb497487",
  1181 => x"dbe4c191",
  1182 => x"c2c1c181",
  1183 => x"ecdcc279",
  1184 => x"d802bf97",
  1185 => x"de497487",
  1186 => x"c284c191",
  1187 => x"714be0e2",
  1188 => x"ecdcc283",
  1189 => x"fe49dd4a",
  1190 => x"d887d5f8",
  1191 => x"de4b7487",
  1192 => x"e0e2c293",
  1193 => x"49a3cb83",
  1194 => x"84c151c0",
  1195 => x"cb4a6e73",
  1196 => x"fbf7fe49",
  1197 => x"4866c487",
  1198 => x"a6c880c1",
  1199 => x"acb7c758",
  1200 => x"87c5c003",
  1201 => x"e2fc056e",
  1202 => x"acb7c787",
  1203 => x"87d9c003",
  1204 => x"48c8e2c2",
  1205 => x"497478c0",
  1206 => x"e2c291de",
  1207 => x"51c081e0",
  1208 => x"b7c784c1",
  1209 => x"e7ff04ac",
  1210 => x"f0e5c187",
  1211 => x"c150c048",
  1212 => x"c148e8e5",
  1213 => x"c178e1cc",
  1214 => x"c148ece5",
  1215 => x"c178e5c2",
  1216 => x"c148f3e5",
  1217 => x"cc78c5c4",
  1218 => x"fbc04966",
  1219 => x"8ef087e2",
  1220 => x"1e87f9e7",
  1221 => x"e1c24a71",
  1222 => x"49725af8",
  1223 => x"2687dbf9",
  1224 => x"4a711e4f",
  1225 => x"c191cb49",
  1226 => x"c881dbe4",
  1227 => x"c2481181",
  1228 => x"c058f4e1",
  1229 => x"fe49a2f0",
  1230 => x"c087c5f6",
  1231 => x"87d5d549",
  1232 => x"5e0e4f26",
  1233 => x"0e5d5c5b",
  1234 => x"4d7186f0",
  1235 => x"c191cb49",
  1236 => x"ca81dbe4",
  1237 => x"a6c47ea1",
  1238 => x"ece1c248",
  1239 => x"976e78bf",
  1240 => x"66c44abf",
  1241 => x"c82b724b",
  1242 => x"48124aa1",
  1243 => x"7058a6cc",
  1244 => x"c983c19b",
  1245 => x"49699781",
  1246 => x"c204abb7",
  1247 => x"6e4bc087",
  1248 => x"c84abf97",
  1249 => x"31724966",
  1250 => x"66c4b9ff",
  1251 => x"724c7399",
  1252 => x"c2b47134",
  1253 => x"ff5cf0e1",
  1254 => x"ffc348d4",
  1255 => x"bfd0ff78",
  1256 => x"c0c0c848",
  1257 => x"58a6d098",
  1258 => x"d0029870",
  1259 => x"bfd0ff87",
  1260 => x"c0c0c848",
  1261 => x"58a6c498",
  1262 => x"f0059870",
  1263 => x"48d0ff87",
  1264 => x"ff78e1c0",
  1265 => x"78de48d4",
  1266 => x"0c7c0c70",
  1267 => x"b7c84874",
  1268 => x"08d4ff28",
  1269 => x"d0487478",
  1270 => x"d4ff28b7",
  1271 => x"48747808",
  1272 => x"ff28b7d8",
  1273 => x"ff7808d4",
  1274 => x"c848bfd0",
  1275 => x"c498c0c0",
  1276 => x"987058a6",
  1277 => x"ff87d002",
  1278 => x"c848bfd0",
  1279 => x"c498c0c0",
  1280 => x"987058a6",
  1281 => x"ff87f005",
  1282 => x"e0c048d0",
  1283 => x"c01ec778",
  1284 => x"dbe4c11e",
  1285 => x"f0e1c21e",
  1286 => x"e9c149bf",
  1287 => x"c0497587",
  1288 => x"e487cdf7",
  1289 => x"87e4e38e",
  1290 => x"711e731e",
  1291 => x"d1fc494b",
  1292 => x"fc497387",
  1293 => x"d7e387cc",
  1294 => x"1e731e87",
  1295 => x"a3c24b71",
  1296 => x"87d6024a",
  1297 => x"c0058ac1",
  1298 => x"e2c287e2",
  1299 => x"db02bfc4",
  1300 => x"88c14887",
  1301 => x"58c8e2c2",
  1302 => x"e2c287d2",
  1303 => x"cb02bfc8",
  1304 => x"c4e2c287",
  1305 => x"80c148bf",
  1306 => x"58c8e2c2",
  1307 => x"1ec01ec7",
  1308 => x"1edbe4c1",
  1309 => x"bff0e1c2",
  1310 => x"7387cb49",
  1311 => x"eff5c049",
  1312 => x"e28ef487",
  1313 => x"5e0e87ca",
  1314 => x"0e5d5c5b",
  1315 => x"dc86d8ff",
  1316 => x"a6c859a6",
  1317 => x"c478c048",
  1318 => x"4d78c080",
  1319 => x"e2c280c4",
  1320 => x"c278bfc4",
  1321 => x"c148c8e2",
  1322 => x"48d4ff78",
  1323 => x"ff78ffc3",
  1324 => x"c848bfd0",
  1325 => x"c498c0c0",
  1326 => x"987058a6",
  1327 => x"ff87d002",
  1328 => x"c848bfd0",
  1329 => x"c498c0c0",
  1330 => x"987058a6",
  1331 => x"ff87f005",
  1332 => x"e1c048d0",
  1333 => x"48d4ff78",
  1334 => x"deff78d4",
  1335 => x"d4ff87e5",
  1336 => x"78ffc348",
  1337 => x"ff48a6d4",
  1338 => x"d478bfd4",
  1339 => x"fbc04866",
  1340 => x"d1c102a8",
  1341 => x"66f8c087",
  1342 => x"6a82c44a",
  1343 => x"c11e727e",
  1344 => x"c448ecc2",
  1345 => x"a1c84966",
  1346 => x"7141204a",
  1347 => x"87f905aa",
  1348 => x"4a265110",
  1349 => x"4866f8c0",
  1350 => x"78d3ccc1",
  1351 => x"81c7496a",
  1352 => x"c15166d4",
  1353 => x"6a1ed81e",
  1354 => x"ff81c849",
  1355 => x"c887ebdd",
  1356 => x"4866d086",
  1357 => x"01a8b7c0",
  1358 => x"4dc187c4",
  1359 => x"66d087c8",
  1360 => x"d488c148",
  1361 => x"66d458a6",
  1362 => x"87e6ca02",
  1363 => x"b766c0c1",
  1364 => x"ddca03ad",
  1365 => x"48d4ff87",
  1366 => x"d478ffc3",
  1367 => x"d4ff48a6",
  1368 => x"66d478bf",
  1369 => x"88c6c148",
  1370 => x"7058a6c4",
  1371 => x"e6c00298",
  1372 => x"88c94887",
  1373 => x"7058a6c4",
  1374 => x"cec40298",
  1375 => x"88c14887",
  1376 => x"7058a6c4",
  1377 => x"e0c10298",
  1378 => x"88c44887",
  1379 => x"987058a6",
  1380 => x"87f7c302",
  1381 => x"d887c5c9",
  1382 => x"c2c10566",
  1383 => x"48d4ff87",
  1384 => x"c078ffc3",
  1385 => x"751eca1e",
  1386 => x"c193cb4b",
  1387 => x"c48366c0",
  1388 => x"496c4ca3",
  1389 => x"87e2dbff",
  1390 => x"1ede1ec1",
  1391 => x"dbff496c",
  1392 => x"86d087d8",
  1393 => x"7bd3ccc1",
  1394 => x"adb766d0",
  1395 => x"c187c504",
  1396 => x"87cfc885",
  1397 => x"c14866d0",
  1398 => x"58a6d488",
  1399 => x"ff87c4c8",
  1400 => x"d887e0da",
  1401 => x"fac758a6",
  1402 => x"e7dcff87",
  1403 => x"58a6cc87",
  1404 => x"a8b766cc",
  1405 => x"cc87c606",
  1406 => x"66c848a6",
  1407 => x"d3dcff78",
  1408 => x"a8ecc087",
  1409 => x"87c3c205",
  1410 => x"c10566d8",
  1411 => x"497587f3",
  1412 => x"f8c091cb",
  1413 => x"a1c48166",
  1414 => x"c84c6a4a",
  1415 => x"66c84aa1",
  1416 => x"e1ccc152",
  1417 => x"48d4ff79",
  1418 => x"d478ffc3",
  1419 => x"d4ff48a6",
  1420 => x"66d478bf",
  1421 => x"87e8c002",
  1422 => x"a8fbc048",
  1423 => x"87e0c002",
  1424 => x"7c9766d4",
  1425 => x"d4ff84c1",
  1426 => x"78ffc348",
  1427 => x"ff48a6d4",
  1428 => x"d478bfd4",
  1429 => x"87c80266",
  1430 => x"a8fbc048",
  1431 => x"87e0ff05",
  1432 => x"c254e0c0",
  1433 => x"97c054c1",
  1434 => x"b766d07c",
  1435 => x"c5c004ad",
  1436 => x"c585c187",
  1437 => x"66d087ed",
  1438 => x"d488c148",
  1439 => x"e2c558a6",
  1440 => x"fed7ff87",
  1441 => x"58a6d887",
  1442 => x"c887d8c5",
  1443 => x"66d84866",
  1444 => x"fdc405a8",
  1445 => x"48a6dc87",
  1446 => x"d9ff78c0",
  1447 => x"a6d887f6",
  1448 => x"efd9ff58",
  1449 => x"a6e4c087",
  1450 => x"a8ecc058",
  1451 => x"87cac005",
  1452 => x"48a6e0c0",
  1453 => x"c07866d4",
  1454 => x"d4ff87c6",
  1455 => x"78ffc348",
  1456 => x"91cb4975",
  1457 => x"4866f8c0",
  1458 => x"a6c48071",
  1459 => x"ca496e58",
  1460 => x"5166d481",
  1461 => x"4966e0c0",
  1462 => x"66d481c1",
  1463 => x"7148c189",
  1464 => x"c1497030",
  1465 => x"c84a6e89",
  1466 => x"97097282",
  1467 => x"e1c20979",
  1468 => x"d449bfec",
  1469 => x"9729b766",
  1470 => x"71484a6a",
  1471 => x"a6e8c098",
  1472 => x"c4486e58",
  1473 => x"58a6c880",
  1474 => x"4cbf66c4",
  1475 => x"c84866d8",
  1476 => x"c002a866",
  1477 => x"e0c087c9",
  1478 => x"78c048a6",
  1479 => x"c087c6c0",
  1480 => x"c148a6e0",
  1481 => x"66e0c078",
  1482 => x"1ee0c01e",
  1483 => x"d5ff4974",
  1484 => x"86c887e8",
  1485 => x"c058a6d8",
  1486 => x"c106a8b7",
  1487 => x"66d487da",
  1488 => x"bf66c484",
  1489 => x"81e0c049",
  1490 => x"c14b8974",
  1491 => x"714af5c2",
  1492 => x"87dce5fe",
  1493 => x"66dc84c2",
  1494 => x"c080c148",
  1495 => x"c058a6e0",
  1496 => x"c14966e4",
  1497 => x"02a97081",
  1498 => x"c087c9c0",
  1499 => x"c048a6e0",
  1500 => x"87c6c078",
  1501 => x"48a6e0c0",
  1502 => x"e0c078c1",
  1503 => x"66c81e66",
  1504 => x"e0c049bf",
  1505 => x"71897481",
  1506 => x"ff49741e",
  1507 => x"c887cbd4",
  1508 => x"a8b7c086",
  1509 => x"87fefe01",
  1510 => x"c00266dc",
  1511 => x"496e87d0",
  1512 => x"66dc81c9",
  1513 => x"c1486e51",
  1514 => x"c078c2cd",
  1515 => x"496e87cc",
  1516 => x"51c281c9",
  1517 => x"d0c1486e",
  1518 => x"66d078e8",
  1519 => x"c004adb7",
  1520 => x"85c187c5",
  1521 => x"d087dcc0",
  1522 => x"88c14866",
  1523 => x"c058a6d4",
  1524 => x"d2ff87d1",
  1525 => x"a6d887ed",
  1526 => x"87c7c058",
  1527 => x"87e3d2ff",
  1528 => x"d458a6d8",
  1529 => x"c9c00266",
  1530 => x"66c0c187",
  1531 => x"f504adb7",
  1532 => x"b7c787e3",
  1533 => x"dfc003ad",
  1534 => x"c8e2c287",
  1535 => x"7578c048",
  1536 => x"c091cb49",
  1537 => x"c48166f8",
  1538 => x"4a6a4aa1",
  1539 => x"c17952c0",
  1540 => x"adb7c785",
  1541 => x"87e1ff04",
  1542 => x"c00266d8",
  1543 => x"f8c087e2",
  1544 => x"cdc14966",
  1545 => x"66f8c081",
  1546 => x"82d5c14a",
  1547 => x"ccc152c0",
  1548 => x"f8c079e1",
  1549 => x"d1c14966",
  1550 => x"f8c2c181",
  1551 => x"87d6c079",
  1552 => x"4966f8c0",
  1553 => x"c081cdc1",
  1554 => x"c14a66f8",
  1555 => x"c2c182d1",
  1556 => x"c9c27aff",
  1557 => x"d0c179d5",
  1558 => x"f8c04af9",
  1559 => x"d8c14966",
  1560 => x"ff797281",
  1561 => x"c848bfd0",
  1562 => x"c498c0c0",
  1563 => x"987058a6",
  1564 => x"87d1c002",
  1565 => x"48bfd0ff",
  1566 => x"98c0c0c8",
  1567 => x"7058a6c4",
  1568 => x"efff0598",
  1569 => x"48d0ff87",
  1570 => x"cc78e0c0",
  1571 => x"d8ff4866",
  1572 => x"f7d1ff8e",
  1573 => x"1ec71e87",
  1574 => x"e4c11ec0",
  1575 => x"e1c21edb",
  1576 => x"ef49bff0",
  1577 => x"e4c187e0",
  1578 => x"e6c049db",
  1579 => x"8ef487d4",
  1580 => x"c91e4f26",
  1581 => x"e2c287fd",
  1582 => x"50c048d0",
  1583 => x"c348d4ff",
  1584 => x"c3c178ff",
  1585 => x"dffe49c6",
  1586 => x"e8fe87c2",
  1587 => x"987087cd",
  1588 => x"fe87cd02",
  1589 => x"7087caf4",
  1590 => x"87c40298",
  1591 => x"87c24ac1",
  1592 => x"9a724ac0",
  1593 => x"c187c802",
  1594 => x"fe49d0c3",
  1595 => x"c287ddde",
  1596 => x"49bfdcd3",
  1597 => x"87e8d5ff",
  1598 => x"48c4e2c2",
  1599 => x"e1c278c0",
  1600 => x"78c048f0",
  1601 => x"87cdfe49",
  1602 => x"c887d4c3",
  1603 => x"e5c087f9",
  1604 => x"f6ff87d2",
  1605 => x"d34f2687",
  1606 => x"42000010",
  1607 => x"a0000010",
  1608 => x"00000028",
  1609 => x"10420000",
  1610 => x"28be0000",
  1611 => x"00000000",
  1612 => x"00104200",
  1613 => x"0028dc00",
  1614 => x"00000000",
  1615 => x"00001042",
  1616 => x"000028fa",
  1617 => x"42000000",
  1618 => x"18000010",
  1619 => x"00000029",
  1620 => x"10420000",
  1621 => x"29360000",
  1622 => x"00000000",
  1623 => x"00104200",
  1624 => x"00295400",
  1625 => x"00000000",
  1626 => x"00001321",
  1627 => x"00000000",
  1628 => x"05000000",
  1629 => x"00000011",
  1630 => x"00000000",
  1631 => x"1e1e0000",
  1632 => x"c487d5c1",
  1633 => x"262658a6",
  1634 => x"4a711e4f",
  1635 => x"c048f0fe",
  1636 => x"7a0acd78",
  1637 => x"dfe6c10a",
  1638 => x"efdbfe49",
  1639 => x"534f2687",
  1640 => x"68207465",
  1641 => x"6c646e61",
  1642 => x"000a7265",
  1643 => x"69206e49",
  1644 => x"7265746e",
  1645 => x"74707572",
  1646 => x"6e6f6320",
  1647 => x"75727473",
  1648 => x"726f7463",
  1649 => x"c11e000a",
  1650 => x"fe49ece6",
  1651 => x"c187fdda",
  1652 => x"fe49fee5",
  1653 => x"4f2687f3",
  1654 => x"bff0fe1e",
  1655 => x"1e4f2648",
  1656 => x"c148f0fe",
  1657 => x"1e4f2678",
  1658 => x"c048f0fe",
  1659 => x"1e4f2678",
  1660 => x"7ac04a71",
  1661 => x"c049a2c4",
  1662 => x"49a2c879",
  1663 => x"a2cc79c0",
  1664 => x"2679c049",
  1665 => x"5b5e0e4f",
  1666 => x"86f80e5c",
  1667 => x"a4c84c71",
  1668 => x"4ba4cc49",
  1669 => x"80c1486b",
  1670 => x"cf58a6c4",
  1671 => x"58a6c898",
  1672 => x"66c44869",
  1673 => x"87d405a8",
  1674 => x"80c1486b",
  1675 => x"cf58a6c4",
  1676 => x"58a6c898",
  1677 => x"66c44869",
  1678 => x"87ec02a8",
  1679 => x"c187e8fe",
  1680 => x"6b49a4d0",
  1681 => x"c490c448",
  1682 => x"817058a6",
  1683 => x"6b7966d4",
  1684 => x"c880c148",
  1685 => x"98cf58a6",
  1686 => x"d2c17b70",
  1687 => x"87fffd87",
  1688 => x"87c28ef8",
  1689 => x"4c264d26",
  1690 => x"4f264b26",
  1691 => x"5c5b5e0e",
  1692 => x"86f80e5d",
  1693 => x"a5c44d71",
  1694 => x"6c486d4c",
  1695 => x"87c505a8",
  1696 => x"e5c048ff",
  1697 => x"87dffd87",
  1698 => x"6c4ba5d0",
  1699 => x"c490c448",
  1700 => x"837058a6",
  1701 => x"ffc34b6b",
  1702 => x"c1486c9b",
  1703 => x"58a6c880",
  1704 => x"7c7098cf",
  1705 => x"7387f8fc",
  1706 => x"8ef84849",
  1707 => x"1e87f5fe",
  1708 => x"86f81e73",
  1709 => x"e087f0fc",
  1710 => x"c0494bbf",
  1711 => x"0299c0e0",
  1712 => x"7387e7c0",
  1713 => x"9affc34a",
  1714 => x"bff2e5c2",
  1715 => x"c490c448",
  1716 => x"e6c258a6",
  1717 => x"817049c2",
  1718 => x"e5c27972",
  1719 => x"c148bff2",
  1720 => x"58a6c880",
  1721 => x"e5c298cf",
  1722 => x"497358f6",
  1723 => x"0299c0d0",
  1724 => x"c287f2c0",
  1725 => x"48bffae5",
  1726 => x"bffee5c2",
  1727 => x"e4c002a8",
  1728 => x"fae5c287",
  1729 => x"90c448bf",
  1730 => x"c258a6c4",
  1731 => x"7049c2e7",
  1732 => x"6948e081",
  1733 => x"fae5c278",
  1734 => x"80c148bf",
  1735 => x"cf58a6c8",
  1736 => x"fee5c298",
  1737 => x"87f0fa58",
  1738 => x"fa58a6c4",
  1739 => x"8ef887f1",
  1740 => x"1e87f5fc",
  1741 => x"49f2e5c2",
  1742 => x"c187f4fa",
  1743 => x"f949efea",
  1744 => x"f5c387c7",
  1745 => x"1e4f2687",
  1746 => x"e5c21e73",
  1747 => x"dbfc49f2",
  1748 => x"c04a7087",
  1749 => x"c204aab7",
  1750 => x"f0c387cc",
  1751 => x"87c905aa",
  1752 => x"48f2efc1",
  1753 => x"edc178c1",
  1754 => x"aae0c387",
  1755 => x"c187c905",
  1756 => x"c148f6ef",
  1757 => x"87dec178",
  1758 => x"bff6efc1",
  1759 => x"c287c602",
  1760 => x"c24ba2c0",
  1761 => x"c14b7287",
  1762 => x"02bff2ef",
  1763 => x"7387e0c0",
  1764 => x"29b7c449",
  1765 => x"faefc191",
  1766 => x"cf4a7381",
  1767 => x"c192c29a",
  1768 => x"70307248",
  1769 => x"72baff4a",
  1770 => x"70986948",
  1771 => x"7387db79",
  1772 => x"29b7c449",
  1773 => x"faefc191",
  1774 => x"cf4a7381",
  1775 => x"c392c29a",
  1776 => x"70307248",
  1777 => x"b069484a",
  1778 => x"efc17970",
  1779 => x"78c048f6",
  1780 => x"48f2efc1",
  1781 => x"e5c278c0",
  1782 => x"cffa49f2",
  1783 => x"c04a7087",
  1784 => x"fd03aab7",
  1785 => x"48c087f4",
  1786 => x"4d2687c4",
  1787 => x"4b264c26",
  1788 => x"00004f26",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"c01e0000",
  1807 => x"c449724a",
  1808 => x"faefc191",
  1809 => x"c179c081",
  1810 => x"aab7d082",
  1811 => x"2687ee04",
  1812 => x"5b5e0e4f",
  1813 => x"710e5d5c",
  1814 => x"87cbf64d",
  1815 => x"b7c44a75",
  1816 => x"efc1922a",
  1817 => x"4c7582fa",
  1818 => x"94c29ccf",
  1819 => x"744b496a",
  1820 => x"c29bc32b",
  1821 => x"70307448",
  1822 => x"74bcff4c",
  1823 => x"70987148",
  1824 => x"87dbf57a",
  1825 => x"e1fd4873",
  1826 => x"ff1e1e87",
  1827 => x"c848bfd0",
  1828 => x"c498c0c0",
  1829 => x"987058a6",
  1830 => x"ff87d002",
  1831 => x"c848bfd0",
  1832 => x"c498c0c0",
  1833 => x"987058a6",
  1834 => x"ff87f005",
  1835 => x"e1c448d0",
  1836 => x"ff487178",
  1837 => x"c87808d4",
  1838 => x"d4ff4866",
  1839 => x"26267808",
  1840 => x"711e1e4f",
  1841 => x"4966c84a",
  1842 => x"fe49721e",
  1843 => x"86c487fb",
  1844 => x"48bfd0ff",
  1845 => x"98c0c0c8",
  1846 => x"7058a6c4",
  1847 => x"87d00298",
  1848 => x"48bfd0ff",
  1849 => x"98c0c0c8",
  1850 => x"7058a6c4",
  1851 => x"87f00598",
  1852 => x"c048d0ff",
  1853 => x"262678e0",
  1854 => x"1e731e4f",
  1855 => x"66c84b71",
  1856 => x"c14a731e",
  1857 => x"fe49a2e0",
  1858 => x"c42687f7",
  1859 => x"264d2687",
  1860 => x"264b264c",
  1861 => x"ff1e1e4f",
  1862 => x"c848bfd0",
  1863 => x"c498c0c0",
  1864 => x"987058a6",
  1865 => x"ff87d002",
  1866 => x"c848bfd0",
  1867 => x"c498c0c0",
  1868 => x"987058a6",
  1869 => x"ff87f005",
  1870 => x"c9c448d0",
  1871 => x"ff487178",
  1872 => x"267808d4",
  1873 => x"1e1e4f26",
  1874 => x"ff494a71",
  1875 => x"d0ff87c7",
  1876 => x"c0c848bf",
  1877 => x"a6c498c0",
  1878 => x"02987058",
  1879 => x"d0ff87d0",
  1880 => x"c0c848bf",
  1881 => x"a6c498c0",
  1882 => x"05987058",
  1883 => x"d0ff87f0",
  1884 => x"2678c848",
  1885 => x"731e4f26",
  1886 => x"4b711e1e",
  1887 => x"bfcee8c2",
  1888 => x"c387c302",
  1889 => x"d0ff87cc",
  1890 => x"c0c848bf",
  1891 => x"a6c498c0",
  1892 => x"02987058",
  1893 => x"d0ff87d0",
  1894 => x"c0c848bf",
  1895 => x"a6c498c0",
  1896 => x"05987058",
  1897 => x"d0ff87f0",
  1898 => x"78c9c448",
  1899 => x"e0c04873",
  1900 => x"08d4ffb0",
  1901 => x"c2e8c278",
  1902 => x"cc78c048",
  1903 => x"87c50266",
  1904 => x"c249ffc3",
  1905 => x"c249c087",
  1906 => x"d059cae8",
  1907 => x"87c60266",
  1908 => x"4ad5d5c5",
  1909 => x"ffcf87c4",
  1910 => x"e8c24aff",
  1911 => x"e8c25ace",
  1912 => x"78c148ce",
  1913 => x"2687c426",
  1914 => x"264c264d",
  1915 => x"0e4f264b",
  1916 => x"5d5c5b5e",
  1917 => x"c24a710e",
  1918 => x"4cbfcae8",
  1919 => x"cb029a72",
  1920 => x"91c84987",
  1921 => x"4bf0f6c1",
  1922 => x"87c48371",
  1923 => x"4bf0fac1",
  1924 => x"49134dc0",
  1925 => x"e8c29974",
  1926 => x"7148bfc6",
  1927 => x"08d4ffb8",
  1928 => x"2cb7c178",
  1929 => x"adb7c885",
  1930 => x"c287e704",
  1931 => x"48bfc2e8",
  1932 => x"e8c280c8",
  1933 => x"eefe58c6",
  1934 => x"1e731e87",
  1935 => x"4a134b71",
  1936 => x"87cb029a",
  1937 => x"e6fe4972",
  1938 => x"9a4a1387",
  1939 => x"fe87f505",
  1940 => x"1e1e87d9",
  1941 => x"bfc2e8c2",
  1942 => x"c2e8c249",
  1943 => x"78a1c148",
  1944 => x"a9b7c0c4",
  1945 => x"ff87db03",
  1946 => x"e8c248d4",
  1947 => x"c278bfc6",
  1948 => x"49bfc2e8",
  1949 => x"48c2e8c2",
  1950 => x"c478a1c1",
  1951 => x"04a9b7c0",
  1952 => x"d0ff87e5",
  1953 => x"c0c848bf",
  1954 => x"a6c498c0",
  1955 => x"02987058",
  1956 => x"d0ff87d0",
  1957 => x"c0c848bf",
  1958 => x"a6c498c0",
  1959 => x"05987058",
  1960 => x"d0ff87f0",
  1961 => x"c278c848",
  1962 => x"c048cee8",
  1963 => x"4f262678",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"5f000000",
  1967 => x"0000005f",
  1968 => x"00030300",
  1969 => x"00000303",
  1970 => x"147f7f14",
  1971 => x"00147f7f",
  1972 => x"6b2e2400",
  1973 => x"00123a6b",
  1974 => x"18366a4c",
  1975 => x"0032566c",
  1976 => x"594f7e30",
  1977 => x"40683a77",
  1978 => x"07040000",
  1979 => x"00000003",
  1980 => x"3e1c0000",
  1981 => x"00004163",
  1982 => x"63410000",
  1983 => x"00001c3e",
  1984 => x"1c3e2a08",
  1985 => x"082a3e1c",
  1986 => x"3e080800",
  1987 => x"0008083e",
  1988 => x"e0800000",
  1989 => x"00000060",
  1990 => x"08080800",
  1991 => x"00080808",
  1992 => x"60000000",
  1993 => x"00000060",
  1994 => x"18306040",
  1995 => x"0103060c",
  1996 => x"597f3e00",
  1997 => x"003e7f4d",
  1998 => x"7f060400",
  1999 => x"0000007f",
  2000 => x"71634200",
  2001 => x"00464f59",
  2002 => x"49632200",
  2003 => x"00367f49",
  2004 => x"13161c18",
  2005 => x"00107f7f",
  2006 => x"45672700",
  2007 => x"00397d45",
  2008 => x"4b7e3c00",
  2009 => x"00307949",
  2010 => x"71010100",
  2011 => x"00070f79",
  2012 => x"497f3600",
  2013 => x"00367f49",
  2014 => x"494f0600",
  2015 => x"001e3f69",
  2016 => x"66000000",
  2017 => x"00000066",
  2018 => x"e6800000",
  2019 => x"00000066",
  2020 => x"14080800",
  2021 => x"00222214",
  2022 => x"14141400",
  2023 => x"00141414",
  2024 => x"14222200",
  2025 => x"00080814",
  2026 => x"51030200",
  2027 => x"00060f59",
  2028 => x"5d417f3e",
  2029 => x"001e1f55",
  2030 => x"097f7e00",
  2031 => x"007e7f09",
  2032 => x"497f7f00",
  2033 => x"00367f49",
  2034 => x"633e1c00",
  2035 => x"00414141",
  2036 => x"417f7f00",
  2037 => x"001c3e63",
  2038 => x"497f7f00",
  2039 => x"00414149",
  2040 => x"097f7f00",
  2041 => x"00010109",
  2042 => x"417f3e00",
  2043 => x"007a7b49",
  2044 => x"087f7f00",
  2045 => x"007f7f08",
  2046 => x"7f410000",
  2047 => x"0000417f",
  2048 => x"40602000",
  2049 => x"003f7f40",
  2050 => x"1c087f7f",
  2051 => x"00416336",
  2052 => x"407f7f00",
  2053 => x"00404040",
  2054 => x"0c067f7f",
  2055 => x"007f7f06",
  2056 => x"0c067f7f",
  2057 => x"007f7f18",
  2058 => x"417f3e00",
  2059 => x"003e7f41",
  2060 => x"097f7f00",
  2061 => x"00060f09",
  2062 => x"61417f3e",
  2063 => x"00407e7f",
  2064 => x"097f7f00",
  2065 => x"00667f19",
  2066 => x"4d6f2600",
  2067 => x"00327b59",
  2068 => x"7f010100",
  2069 => x"0001017f",
  2070 => x"407f3f00",
  2071 => x"003f7f40",
  2072 => x"703f0f00",
  2073 => x"000f3f70",
  2074 => x"18307f7f",
  2075 => x"007f7f30",
  2076 => x"1c366341",
  2077 => x"4163361c",
  2078 => x"7c060301",
  2079 => x"0103067c",
  2080 => x"4d597161",
  2081 => x"00414347",
  2082 => x"7f7f0000",
  2083 => x"00004141",
  2084 => x"0c060301",
  2085 => x"40603018",
  2086 => x"41410000",
  2087 => x"00007f7f",
  2088 => x"03060c08",
  2089 => x"00080c06",
  2090 => x"80808080",
  2091 => x"00808080",
  2092 => x"03000000",
  2093 => x"00000407",
  2094 => x"54742000",
  2095 => x"00787c54",
  2096 => x"447f7f00",
  2097 => x"00387c44",
  2098 => x"447c3800",
  2099 => x"00004444",
  2100 => x"447c3800",
  2101 => x"007f7f44",
  2102 => x"547c3800",
  2103 => x"00185c54",
  2104 => x"7f7e0400",
  2105 => x"00000505",
  2106 => x"a4bc1800",
  2107 => x"007cfca4",
  2108 => x"047f7f00",
  2109 => x"00787c04",
  2110 => x"3d000000",
  2111 => x"0000407d",
  2112 => x"80808000",
  2113 => x"00007dfd",
  2114 => x"107f7f00",
  2115 => x"00446c38",
  2116 => x"3f000000",
  2117 => x"0000407f",
  2118 => x"180c7c7c",
  2119 => x"00787c0c",
  2120 => x"047c7c00",
  2121 => x"00787c04",
  2122 => x"447c3800",
  2123 => x"00387c44",
  2124 => x"24fcfc00",
  2125 => x"00183c24",
  2126 => x"243c1800",
  2127 => x"00fcfc24",
  2128 => x"047c7c00",
  2129 => x"00080c04",
  2130 => x"545c4800",
  2131 => x"00207454",
  2132 => x"7f3f0400",
  2133 => x"00004444",
  2134 => x"407c3c00",
  2135 => x"007c7c40",
  2136 => x"603c1c00",
  2137 => x"001c3c60",
  2138 => x"30607c3c",
  2139 => x"003c7c60",
  2140 => x"10386c44",
  2141 => x"00446c38",
  2142 => x"e0bc1c00",
  2143 => x"001c3c60",
  2144 => x"74644400",
  2145 => x"00444c5c",
  2146 => x"3e080800",
  2147 => x"00414177",
  2148 => x"7f000000",
  2149 => x"0000007f",
  2150 => x"77414100",
  2151 => x"0008083e",
  2152 => x"03010102",
  2153 => x"00010202",
  2154 => x"7f7f7f7f",
  2155 => x"007f7f7f",
  2156 => x"1c1c0808",
  2157 => x"7f7f3e3e",
  2158 => x"3e3e7f7f",
  2159 => x"08081c1c",
  2160 => x"7c181000",
  2161 => x"0010187c",
  2162 => x"7c301000",
  2163 => x"0010307c",
  2164 => x"60603010",
  2165 => x"00061e78",
  2166 => x"183c6642",
  2167 => x"0042663c",
  2168 => x"c26a3878",
  2169 => x"00386cc6",
  2170 => x"60000060",
  2171 => x"00600000",
  2172 => x"5c5b5e0e",
  2173 => x"711e0e5d",
  2174 => x"d6e8c24c",
  2175 => x"4bc04dbf",
  2176 => x"ab741ec0",
  2177 => x"c487c702",
  2178 => x"78c048a6",
  2179 => x"a6c487c5",
  2180 => x"c478c148",
  2181 => x"49731e66",
  2182 => x"c887dbed",
  2183 => x"49e0c086",
  2184 => x"c487ccef",
  2185 => x"496a4aa5",
  2186 => x"f087cef0",
  2187 => x"85cb87e4",
  2188 => x"b7c883c1",
  2189 => x"c7ff04ab",
  2190 => x"4d262687",
  2191 => x"4b264c26",
  2192 => x"711e4f26",
  2193 => x"dae8c24a",
  2194 => x"dae8c25a",
  2195 => x"4978c748",
  2196 => x"2687ddfe",
  2197 => x"c0c11e4f",
  2198 => x"87eaeb49",
  2199 => x"48c5d3c2",
  2200 => x"4f2678c0",
  2201 => x"5c5b5e0e",
  2202 => x"86f40e5d",
  2203 => x"a6c87ec0",
  2204 => x"78bfec48",
  2205 => x"e8c280fc",
  2206 => x"c278bfd6",
  2207 => x"4dbfdee8",
  2208 => x"c74cbfe8",
  2209 => x"87c9e749",
  2210 => x"99c24970",
  2211 => x"c287d005",
  2212 => x"49bffdd2",
  2213 => x"66c8b9ff",
  2214 => x"0299c199",
  2215 => x"c787ebc0",
  2216 => x"87ede649",
  2217 => x"cd029870",
  2218 => x"87dbe287",
  2219 => x"e0e649c7",
  2220 => x"05987087",
  2221 => x"d3c287f3",
  2222 => x"c14abfc5",
  2223 => x"c9d3c2ba",
  2224 => x"a2c0c15a",
  2225 => x"87fee949",
  2226 => x"d2c27ec1",
  2227 => x"66c848fd",
  2228 => x"c5d3c278",
  2229 => x"cbc105bf",
  2230 => x"c0c0c887",
  2231 => x"c9d3c27e",
  2232 => x"e549134b",
  2233 => x"987087eb",
  2234 => x"6e87c202",
  2235 => x"c1486eb4",
  2236 => x"a6c428b7",
  2237 => x"05987058",
  2238 => x"7487e6ff",
  2239 => x"99ffc349",
  2240 => x"49c01e71",
  2241 => x"7487f2e7",
  2242 => x"29b7c849",
  2243 => x"49c11e71",
  2244 => x"c887e6e7",
  2245 => x"49fdc386",
  2246 => x"c387f6e4",
  2247 => x"f0e449fa",
  2248 => x"87c4c687",
  2249 => x"ffc34974",
  2250 => x"2cb7c899",
  2251 => x"9c74b471",
  2252 => x"87e2c002",
  2253 => x"ff48a6c8",
  2254 => x"c878bfc8",
  2255 => x"d3c24966",
  2256 => x"c289bfc1",
  2257 => x"c403a9e0",
  2258 => x"cf4cc087",
  2259 => x"c1d3c287",
  2260 => x"7866c848",
  2261 => x"d3c287c6",
  2262 => x"78c048c1",
  2263 => x"99c84974",
  2264 => x"c387ce05",
  2265 => x"e8e349f5",
  2266 => x"c2497087",
  2267 => x"e6c00299",
  2268 => x"dae8c287",
  2269 => x"87c902bf",
  2270 => x"c288c148",
  2271 => x"d458dee8",
  2272 => x"4866c487",
  2273 => x"c480d8c1",
  2274 => x"bf6e58a6",
  2275 => x"87c5c002",
  2276 => x"7349ff4b",
  2277 => x"747ec10f",
  2278 => x"0599c449",
  2279 => x"f2c387ce",
  2280 => x"87ede249",
  2281 => x"99c24970",
  2282 => x"87eec002",
  2283 => x"bfdae8c2",
  2284 => x"c7486e7e",
  2285 => x"c003a8b7",
  2286 => x"486e87ca",
  2287 => x"e8c280c1",
  2288 => x"87d458de",
  2289 => x"c14866c4",
  2290 => x"a6c480d8",
  2291 => x"02bf6e58",
  2292 => x"4b87c5c0",
  2293 => x"0f7349fe",
  2294 => x"fdc37ec1",
  2295 => x"87f1e149",
  2296 => x"99c24970",
  2297 => x"87e3c002",
  2298 => x"bfdae8c2",
  2299 => x"87c9c002",
  2300 => x"48dae8c2",
  2301 => x"d0c078c0",
  2302 => x"4a66c487",
  2303 => x"6a82d8c1",
  2304 => x"87c5c002",
  2305 => x"7349fd4b",
  2306 => x"c37ec10f",
  2307 => x"c0e149fa",
  2308 => x"c2497087",
  2309 => x"ebc00299",
  2310 => x"dae8c287",
  2311 => x"b7c748bf",
  2312 => x"c9c003a8",
  2313 => x"dae8c287",
  2314 => x"c078c748",
  2315 => x"66c487d4",
  2316 => x"80d8c148",
  2317 => x"6e58a6c4",
  2318 => x"c5c002bf",
  2319 => x"49fc4b87",
  2320 => x"7ec10f73",
  2321 => x"f0c34974",
  2322 => x"cfc00599",
  2323 => x"49dac187",
  2324 => x"87fddfff",
  2325 => x"99c24970",
  2326 => x"87d0c002",
  2327 => x"bfdae8c2",
  2328 => x"93cb4b49",
  2329 => x"6b8366c4",
  2330 => x"0f73714b",
  2331 => x"c0029d75",
  2332 => x"026d87e9",
  2333 => x"6d87e4c0",
  2334 => x"d4dfff49",
  2335 => x"c1497087",
  2336 => x"cbc00299",
  2337 => x"4ba5c487",
  2338 => x"bfdae8c2",
  2339 => x"0f4b6b49",
  2340 => x"c00285c8",
  2341 => x"056d87c5",
  2342 => x"6e87dcff",
  2343 => x"87c8c002",
  2344 => x"bfdae8c2",
  2345 => x"87c8f549",
  2346 => x"cdf68ef4",
  2347 => x"11125887",
  2348 => x"1c1b1d14",
  2349 => x"91595a23",
  2350 => x"ebf2f594",
  2351 => x"000000f4",
  2352 => x"00000000",
  2353 => x"00000000",
  2354 => x"14125800",
  2355 => x"1c1b1d11",
  2356 => x"94595a23",
  2357 => x"ebf2f591",
  2358 => x"000000f4",
  2359 => x"000024e0",
  2360 => x"4f545541",
  2361 => x"544f4f42",
  2362 => x"0053454e",
  2363 => x"000019c6",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
