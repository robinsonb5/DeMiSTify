../demistify_config_pkg.vhd