
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e4",x"e8",x"c2",x"87"),
    12 => (x"48",x"c0",x"c4",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"05",x"88"),
    17 => (x"49",x"e4",x"e8",x"c2"),
    18 => (x"48",x"f0",x"d3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"f0",x"d3",x"c2",x"87"),
    25 => (x"ec",x"d3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e0",x"c1",x"87",x"f7"),
    29 => (x"d3",x"c2",x"87",x"fc"),
    30 => (x"d3",x"c2",x"4d",x"f0"),
    31 => (x"ad",x"74",x"4c",x"f0"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"c0",x"4b",x"71",x"0e"),
    37 => (x"9a",x"4a",x"13",x"4c"),
    38 => (x"72",x"87",x"cd",x"02"),
    39 => (x"87",x"e0",x"c0",x"49"),
    40 => (x"4a",x"13",x"84",x"c1"),
    41 => (x"87",x"f3",x"05",x"9a"),
    42 => (x"4c",x"26",x"48",x"74"),
    43 => (x"4f",x"26",x"4b",x"26"),
    44 => (x"81",x"48",x"73",x"1e"),
    45 => (x"c5",x"02",x"a9",x"73"),
    46 => (x"05",x"53",x"12",x"87"),
    47 => (x"4f",x"26",x"87",x"f6"),
    48 => (x"c0",x"ff",x"1e",x"1e"),
    49 => (x"c4",x"48",x"6a",x"4a"),
    50 => (x"a6",x"c4",x"98",x"c0"),
    51 => (x"02",x"98",x"70",x"58"),
    52 => (x"7a",x"71",x"87",x"f3"),
    53 => (x"4f",x"26",x"26",x"48"),
    54 => (x"ff",x"1e",x"73",x"1e"),
    55 => (x"ff",x"c3",x"4b",x"d4"),
    56 => (x"c3",x"4a",x"6b",x"7b"),
    57 => (x"49",x"6b",x"7b",x"ff"),
    58 => (x"b1",x"72",x"32",x"c8"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"71",x"31",x"c8",x"4a"),
    61 => (x"7b",x"ff",x"c3",x"b2"),
    62 => (x"32",x"c8",x"49",x"6b"),
    63 => (x"48",x"71",x"b1",x"72"),
    64 => (x"4d",x"26",x"87",x"c4"),
    65 => (x"4b",x"26",x"4c",x"26"),
    66 => (x"5e",x"0e",x"4f",x"26"),
    67 => (x"0e",x"5d",x"5c",x"5b"),
    68 => (x"d4",x"ff",x"4a",x"71"),
    69 => (x"c3",x"48",x"72",x"4c"),
    70 => (x"7c",x"70",x"98",x"ff"),
    71 => (x"bf",x"f0",x"d3",x"c2"),
    72 => (x"d0",x"87",x"c8",x"05"),
    73 => (x"30",x"c9",x"48",x"66"),
    74 => (x"d0",x"58",x"a6",x"d4"),
    75 => (x"29",x"d8",x"49",x"66"),
    76 => (x"ff",x"c3",x"48",x"71"),
    77 => (x"d0",x"7c",x"70",x"98"),
    78 => (x"29",x"d0",x"49",x"66"),
    79 => (x"ff",x"c3",x"48",x"71"),
    80 => (x"d0",x"7c",x"70",x"98"),
    81 => (x"29",x"c8",x"49",x"66"),
    82 => (x"ff",x"c3",x"48",x"71"),
    83 => (x"d0",x"7c",x"70",x"98"),
    84 => (x"ff",x"c3",x"48",x"66"),
    85 => (x"72",x"7c",x"70",x"98"),
    86 => (x"71",x"29",x"d0",x"49"),
    87 => (x"98",x"ff",x"c3",x"48"),
    88 => (x"4b",x"6c",x"7c",x"70"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"ff",x"fd"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"df",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c1",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"de",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"49",x"e3",x"c8",x"78"),
   125 => (x"d3",x"87",x"d5",x"fa"),
   126 => (x"c0",x"1e",x"c0",x"4b"),
   127 => (x"c1",x"c1",x"f0",x"ff"),
   128 => (x"87",x"c6",x"fc",x"49"),
   129 => (x"98",x"70",x"86",x"c4"),
   130 => (x"ff",x"87",x"ca",x"05"),
   131 => (x"ff",x"c3",x"48",x"d4"),
   132 => (x"cb",x"48",x"c1",x"78"),
   133 => (x"87",x"eb",x"fd",x"87"),
   134 => (x"ff",x"05",x"8b",x"c1"),
   135 => (x"48",x"c0",x"87",x"db"),
   136 => (x"43",x"87",x"e3",x"fb"),
   137 => (x"53",x"00",x"44",x"4d"),
   138 => (x"20",x"43",x"48",x"44"),
   139 => (x"6c",x"69",x"61",x"66"),
   140 => (x"49",x"00",x"0a",x"21"),
   141 => (x"00",x"52",x"52",x"45"),
   142 => (x"00",x"49",x"50",x"53"),
   143 => (x"74",x"69",x"72",x"57"),
   144 => (x"61",x"66",x"20",x"65"),
   145 => (x"64",x"65",x"6c",x"69"),
   146 => (x"5e",x"0e",x"00",x"0a"),
   147 => (x"ff",x"0e",x"5c",x"5b"),
   148 => (x"ee",x"fc",x"4c",x"d4"),
   149 => (x"1e",x"ea",x"c6",x"87"),
   150 => (x"c1",x"f0",x"e1",x"c0"),
   151 => (x"e9",x"fa",x"49",x"c8"),
   152 => (x"c1",x"86",x"c4",x"87"),
   153 => (x"87",x"c8",x"02",x"a8"),
   154 => (x"c0",x"87",x"fd",x"fd"),
   155 => (x"87",x"e8",x"c1",x"48"),
   156 => (x"70",x"87",x"e5",x"f9"),
   157 => (x"ff",x"ff",x"cf",x"49"),
   158 => (x"a9",x"ea",x"c6",x"99"),
   159 => (x"fd",x"87",x"c8",x"02"),
   160 => (x"48",x"c0",x"87",x"e6"),
   161 => (x"c3",x"87",x"d1",x"c1"),
   162 => (x"f1",x"c0",x"7c",x"ff"),
   163 => (x"87",x"c7",x"fc",x"4b"),
   164 => (x"c0",x"02",x"98",x"70"),
   165 => (x"1e",x"c0",x"87",x"eb"),
   166 => (x"c1",x"f0",x"ff",x"c0"),
   167 => (x"e9",x"f9",x"49",x"fa"),
   168 => (x"70",x"86",x"c4",x"87"),
   169 => (x"87",x"d9",x"05",x"98"),
   170 => (x"6c",x"7c",x"ff",x"c3"),
   171 => (x"7c",x"ff",x"c3",x"49"),
   172 => (x"c1",x"7c",x"7c",x"7c"),
   173 => (x"c4",x"02",x"99",x"c0"),
   174 => (x"db",x"48",x"c1",x"87"),
   175 => (x"d7",x"48",x"c0",x"87"),
   176 => (x"05",x"ab",x"c2",x"87"),
   177 => (x"e7",x"c8",x"87",x"ca"),
   178 => (x"87",x"c0",x"f7",x"49"),
   179 => (x"87",x"c8",x"48",x"c0"),
   180 => (x"fe",x"05",x"8b",x"c1"),
   181 => (x"48",x"c0",x"87",x"f7"),
   182 => (x"0e",x"87",x"e9",x"f8"),
   183 => (x"5d",x"5c",x"5b",x"5e"),
   184 => (x"d0",x"ff",x"1e",x"0e"),
   185 => (x"c0",x"c0",x"c8",x"4d"),
   186 => (x"f0",x"d3",x"c2",x"4b"),
   187 => (x"c8",x"78",x"c1",x"48"),
   188 => (x"d7",x"f6",x"49",x"f8"),
   189 => (x"6d",x"4c",x"c7",x"87"),
   190 => (x"c4",x"98",x"73",x"48"),
   191 => (x"98",x"70",x"58",x"a6"),
   192 => (x"6d",x"87",x"cc",x"02"),
   193 => (x"c4",x"98",x"73",x"48"),
   194 => (x"98",x"70",x"58",x"a6"),
   195 => (x"c2",x"87",x"f4",x"05"),
   196 => (x"87",x"ef",x"f9",x"7d"),
   197 => (x"98",x"73",x"48",x"6d"),
   198 => (x"70",x"58",x"a6",x"c4"),
   199 => (x"87",x"cc",x"02",x"98"),
   200 => (x"98",x"73",x"48",x"6d"),
   201 => (x"70",x"58",x"a6",x"c4"),
   202 => (x"87",x"f4",x"05",x"98"),
   203 => (x"1e",x"c0",x"7d",x"c3"),
   204 => (x"c1",x"d0",x"e5",x"c0"),
   205 => (x"d1",x"f7",x"49",x"c0"),
   206 => (x"c1",x"86",x"c4",x"87"),
   207 => (x"87",x"c1",x"05",x"a8"),
   208 => (x"05",x"ac",x"c2",x"4c"),
   209 => (x"f3",x"c8",x"87",x"cb"),
   210 => (x"87",x"c0",x"f5",x"49"),
   211 => (x"ce",x"c1",x"48",x"c0"),
   212 => (x"05",x"8c",x"c1",x"87"),
   213 => (x"fb",x"87",x"e0",x"fe"),
   214 => (x"d3",x"c2",x"87",x"f0"),
   215 => (x"98",x"70",x"58",x"f4"),
   216 => (x"c1",x"87",x"cd",x"05"),
   217 => (x"f0",x"ff",x"c0",x"1e"),
   218 => (x"f6",x"49",x"d0",x"c1"),
   219 => (x"86",x"c4",x"87",x"dc"),
   220 => (x"c3",x"48",x"d4",x"ff"),
   221 => (x"dd",x"c5",x"78",x"ff"),
   222 => (x"f8",x"d3",x"c2",x"87"),
   223 => (x"73",x"48",x"6d",x"58"),
   224 => (x"58",x"a6",x"c4",x"98"),
   225 => (x"cc",x"02",x"98",x"70"),
   226 => (x"73",x"48",x"6d",x"87"),
   227 => (x"58",x"a6",x"c4",x"98"),
   228 => (x"f4",x"05",x"98",x"70"),
   229 => (x"ff",x"7d",x"c2",x"87"),
   230 => (x"ff",x"c3",x"48",x"d4"),
   231 => (x"26",x"48",x"c1",x"78"),
   232 => (x"0e",x"87",x"df",x"f5"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"c8",x"1e",x"0e"),
   235 => (x"4c",x"c0",x"4b",x"c0"),
   236 => (x"df",x"cd",x"ee",x"c5"),
   237 => (x"5c",x"a6",x"c4",x"4a"),
   238 => (x"c3",x"4c",x"d4",x"ff"),
   239 => (x"48",x"6c",x"7c",x"ff"),
   240 => (x"05",x"a8",x"fe",x"c3"),
   241 => (x"71",x"87",x"c0",x"c2"),
   242 => (x"e2",x"c0",x"05",x"99"),
   243 => (x"bf",x"d0",x"ff",x"87"),
   244 => (x"c4",x"98",x"73",x"48"),
   245 => (x"98",x"70",x"58",x"a6"),
   246 => (x"ff",x"87",x"ce",x"02"),
   247 => (x"73",x"48",x"bf",x"d0"),
   248 => (x"58",x"a6",x"c4",x"98"),
   249 => (x"f2",x"05",x"98",x"70"),
   250 => (x"48",x"d0",x"ff",x"87"),
   251 => (x"d4",x"78",x"d1",x"c4"),
   252 => (x"b7",x"c0",x"48",x"66"),
   253 => (x"e0",x"c0",x"06",x"a8"),
   254 => (x"7c",x"ff",x"c3",x"87"),
   255 => (x"99",x"71",x"4a",x"6c"),
   256 => (x"71",x"87",x"c7",x"02"),
   257 => (x"0a",x"7a",x"97",x"0a"),
   258 => (x"66",x"d4",x"81",x"c1"),
   259 => (x"d8",x"88",x"c1",x"48"),
   260 => (x"b7",x"c0",x"58",x"a6"),
   261 => (x"e0",x"ff",x"01",x"a8"),
   262 => (x"7c",x"ff",x"c3",x"87"),
   263 => (x"05",x"99",x"71",x"7c"),
   264 => (x"ff",x"87",x"e1",x"c0"),
   265 => (x"73",x"48",x"bf",x"d0"),
   266 => (x"58",x"a6",x"c4",x"98"),
   267 => (x"ce",x"02",x"98",x"70"),
   268 => (x"bf",x"d0",x"ff",x"87"),
   269 => (x"c4",x"98",x"73",x"48"),
   270 => (x"98",x"70",x"58",x"a6"),
   271 => (x"ff",x"87",x"f2",x"05"),
   272 => (x"78",x"d0",x"48",x"d0"),
   273 => (x"c1",x"7e",x"4a",x"c1"),
   274 => (x"ee",x"fd",x"05",x"8a"),
   275 => (x"26",x"48",x"6e",x"87"),
   276 => (x"0e",x"87",x"ef",x"f2"),
   277 => (x"0e",x"5c",x"5b",x"5e"),
   278 => (x"c8",x"4a",x"71",x"1e"),
   279 => (x"c0",x"4b",x"c0",x"c0"),
   280 => (x"48",x"d4",x"ff",x"4c"),
   281 => (x"ff",x"78",x"ff",x"c3"),
   282 => (x"73",x"48",x"bf",x"d0"),
   283 => (x"58",x"a6",x"c4",x"98"),
   284 => (x"ce",x"02",x"98",x"70"),
   285 => (x"bf",x"d0",x"ff",x"87"),
   286 => (x"c4",x"98",x"73",x"48"),
   287 => (x"98",x"70",x"58",x"a6"),
   288 => (x"ff",x"87",x"f2",x"05"),
   289 => (x"c3",x"c4",x"48",x"d0"),
   290 => (x"48",x"d4",x"ff",x"78"),
   291 => (x"72",x"78",x"ff",x"c3"),
   292 => (x"f0",x"ff",x"c0",x"1e"),
   293 => (x"f1",x"49",x"d1",x"c1"),
   294 => (x"86",x"c4",x"87",x"f0"),
   295 => (x"c0",x"05",x"98",x"70"),
   296 => (x"c0",x"c8",x"87",x"ee"),
   297 => (x"49",x"66",x"d4",x"1e"),
   298 => (x"c4",x"87",x"f8",x"fb"),
   299 => (x"ff",x"4c",x"70",x"86"),
   300 => (x"73",x"48",x"bf",x"d0"),
   301 => (x"58",x"a6",x"c4",x"98"),
   302 => (x"ce",x"02",x"98",x"70"),
   303 => (x"bf",x"d0",x"ff",x"87"),
   304 => (x"c4",x"98",x"73",x"48"),
   305 => (x"98",x"70",x"58",x"a6"),
   306 => (x"ff",x"87",x"f2",x"05"),
   307 => (x"78",x"c2",x"48",x"d0"),
   308 => (x"f0",x"26",x"48",x"74"),
   309 => (x"5e",x"0e",x"87",x"ee"),
   310 => (x"0e",x"5d",x"5c",x"5b"),
   311 => (x"ff",x"c0",x"1e",x"c0"),
   312 => (x"49",x"c9",x"c1",x"f0"),
   313 => (x"d2",x"87",x"e3",x"f0"),
   314 => (x"fe",x"d3",x"c2",x"1e"),
   315 => (x"87",x"f3",x"fa",x"49"),
   316 => (x"4c",x"c0",x"86",x"c8"),
   317 => (x"b7",x"d2",x"84",x"c1"),
   318 => (x"87",x"f8",x"04",x"ac"),
   319 => (x"97",x"fe",x"d3",x"c2"),
   320 => (x"c0",x"c3",x"49",x"bf"),
   321 => (x"a9",x"c0",x"c1",x"99"),
   322 => (x"87",x"e7",x"c0",x"05"),
   323 => (x"97",x"c5",x"d4",x"c2"),
   324 => (x"31",x"d0",x"49",x"bf"),
   325 => (x"97",x"c6",x"d4",x"c2"),
   326 => (x"32",x"c8",x"4a",x"bf"),
   327 => (x"d4",x"c2",x"b1",x"72"),
   328 => (x"4a",x"bf",x"97",x"c7"),
   329 => (x"cf",x"4c",x"71",x"b1"),
   330 => (x"9c",x"ff",x"ff",x"ff"),
   331 => (x"34",x"ca",x"84",x"c1"),
   332 => (x"c2",x"87",x"e7",x"c1"),
   333 => (x"bf",x"97",x"c7",x"d4"),
   334 => (x"c6",x"31",x"c1",x"49"),
   335 => (x"c8",x"d4",x"c2",x"99"),
   336 => (x"c7",x"4a",x"bf",x"97"),
   337 => (x"b1",x"72",x"2a",x"b7"),
   338 => (x"97",x"c3",x"d4",x"c2"),
   339 => (x"cf",x"4d",x"4a",x"bf"),
   340 => (x"c4",x"d4",x"c2",x"9d"),
   341 => (x"c3",x"4a",x"bf",x"97"),
   342 => (x"c2",x"32",x"ca",x"9a"),
   343 => (x"bf",x"97",x"c5",x"d4"),
   344 => (x"73",x"33",x"c2",x"4b"),
   345 => (x"c6",x"d4",x"c2",x"b2"),
   346 => (x"c3",x"4b",x"bf",x"97"),
   347 => (x"b7",x"c6",x"9b",x"c0"),
   348 => (x"c2",x"b2",x"73",x"2b"),
   349 => (x"71",x"48",x"c1",x"81"),
   350 => (x"c1",x"49",x"70",x"30"),
   351 => (x"70",x"30",x"75",x"48"),
   352 => (x"c1",x"4c",x"72",x"4d"),
   353 => (x"c8",x"94",x"71",x"84"),
   354 => (x"06",x"ad",x"b7",x"c0"),
   355 => (x"34",x"c1",x"87",x"cc"),
   356 => (x"c0",x"c8",x"2d",x"b7"),
   357 => (x"ff",x"01",x"ad",x"b7"),
   358 => (x"48",x"74",x"87",x"f4"),
   359 => (x"0e",x"87",x"e3",x"ed"),
   360 => (x"0e",x"5c",x"5b",x"5e"),
   361 => (x"4c",x"c0",x"4b",x"71"),
   362 => (x"c0",x"48",x"66",x"d0"),
   363 => (x"c0",x"06",x"a8",x"b7"),
   364 => (x"4a",x"13",x"87",x"e3"),
   365 => (x"bf",x"97",x"66",x"cc"),
   366 => (x"48",x"66",x"cc",x"49"),
   367 => (x"a6",x"d0",x"80",x"c1"),
   368 => (x"aa",x"b7",x"71",x"58"),
   369 => (x"c1",x"87",x"c4",x"02"),
   370 => (x"c1",x"87",x"cc",x"48"),
   371 => (x"b7",x"66",x"d0",x"84"),
   372 => (x"dd",x"ff",x"04",x"ac"),
   373 => (x"c2",x"48",x"c0",x"87"),
   374 => (x"26",x"4d",x"26",x"87"),
   375 => (x"26",x"4b",x"26",x"4c"),
   376 => (x"5b",x"5e",x"0e",x"4f"),
   377 => (x"c2",x"0e",x"5d",x"5c"),
   378 => (x"c0",x"48",x"e4",x"dc"),
   379 => (x"dc",x"d4",x"c2",x"78"),
   380 => (x"f9",x"49",x"c0",x"1e"),
   381 => (x"86",x"c4",x"87",x"dd"),
   382 => (x"c5",x"05",x"98",x"70"),
   383 => (x"c8",x"48",x"c0",x"87"),
   384 => (x"4b",x"c0",x"87",x"ef"),
   385 => (x"48",x"dc",x"e1",x"c2"),
   386 => (x"1e",x"c8",x"78",x"c1"),
   387 => (x"1e",x"fd",x"e0",x"c0"),
   388 => (x"49",x"d2",x"d5",x"c2"),
   389 => (x"c8",x"87",x"c8",x"fe"),
   390 => (x"05",x"98",x"70",x"86"),
   391 => (x"e1",x"c2",x"87",x"c6"),
   392 => (x"78",x"c0",x"48",x"dc"),
   393 => (x"e1",x"c0",x"1e",x"c8"),
   394 => (x"d5",x"c2",x"1e",x"c6"),
   395 => (x"ee",x"fd",x"49",x"ee"),
   396 => (x"70",x"86",x"c8",x"87"),
   397 => (x"87",x"c6",x"05",x"98"),
   398 => (x"48",x"dc",x"e1",x"c2"),
   399 => (x"e1",x"c2",x"78",x"c0"),
   400 => (x"c0",x"02",x"bf",x"dc"),
   401 => (x"db",x"c2",x"87",x"fa"),
   402 => (x"c2",x"4b",x"bf",x"e2"),
   403 => (x"bf",x"9f",x"da",x"dc"),
   404 => (x"ea",x"d6",x"c5",x"4a"),
   405 => (x"87",x"c7",x"05",x"aa"),
   406 => (x"bf",x"e2",x"db",x"c2"),
   407 => (x"ca",x"87",x"cc",x"4b"),
   408 => (x"02",x"aa",x"d5",x"e9"),
   409 => (x"48",x"c0",x"87",x"c5"),
   410 => (x"c2",x"87",x"c6",x"c7"),
   411 => (x"73",x"1e",x"dc",x"d4"),
   412 => (x"87",x"df",x"f7",x"49"),
   413 => (x"98",x"70",x"86",x"c4"),
   414 => (x"c0",x"87",x"c5",x"05"),
   415 => (x"87",x"f1",x"c6",x"48"),
   416 => (x"e1",x"c0",x"1e",x"c8"),
   417 => (x"d5",x"c2",x"1e",x"cf"),
   418 => (x"d2",x"fc",x"49",x"ee"),
   419 => (x"70",x"86",x"c8",x"87"),
   420 => (x"87",x"c8",x"05",x"98"),
   421 => (x"48",x"e4",x"dc",x"c2"),
   422 => (x"87",x"da",x"78",x"c1"),
   423 => (x"e1",x"c0",x"1e",x"c8"),
   424 => (x"d5",x"c2",x"1e",x"d8"),
   425 => (x"f6",x"fb",x"49",x"d2"),
   426 => (x"70",x"86",x"c8",x"87"),
   427 => (x"c5",x"c0",x"02",x"98"),
   428 => (x"c5",x"48",x"c0",x"87"),
   429 => (x"dc",x"c2",x"87",x"fb"),
   430 => (x"49",x"bf",x"97",x"da"),
   431 => (x"05",x"a9",x"d5",x"c1"),
   432 => (x"c2",x"87",x"cd",x"c0"),
   433 => (x"bf",x"97",x"db",x"dc"),
   434 => (x"a9",x"ea",x"c2",x"49"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dc",x"c5",x"48",x"c0"),
   437 => (x"dc",x"d4",x"c2",x"87"),
   438 => (x"c3",x"4c",x"bf",x"97"),
   439 => (x"c0",x"02",x"ac",x"e9"),
   440 => (x"eb",x"c3",x"87",x"cc"),
   441 => (x"c5",x"c0",x"02",x"ac"),
   442 => (x"c5",x"48",x"c0",x"87"),
   443 => (x"d4",x"c2",x"87",x"c3"),
   444 => (x"49",x"bf",x"97",x"e7"),
   445 => (x"cc",x"c0",x"05",x"99"),
   446 => (x"e8",x"d4",x"c2",x"87"),
   447 => (x"c2",x"49",x"bf",x"97"),
   448 => (x"c5",x"c0",x"02",x"a9"),
   449 => (x"c4",x"48",x"c0",x"87"),
   450 => (x"d4",x"c2",x"87",x"e7"),
   451 => (x"48",x"bf",x"97",x"e9"),
   452 => (x"58",x"e0",x"dc",x"c2"),
   453 => (x"dc",x"c2",x"88",x"c1"),
   454 => (x"d4",x"c2",x"58",x"e4"),
   455 => (x"49",x"bf",x"97",x"ea"),
   456 => (x"d4",x"c2",x"81",x"73"),
   457 => (x"4a",x"bf",x"97",x"eb"),
   458 => (x"71",x"35",x"c8",x"4d"),
   459 => (x"fc",x"e0",x"c2",x"85"),
   460 => (x"ec",x"d4",x"c2",x"5d"),
   461 => (x"c2",x"48",x"bf",x"97"),
   462 => (x"c2",x"58",x"d0",x"e1"),
   463 => (x"02",x"bf",x"e4",x"dc"),
   464 => (x"c8",x"87",x"dc",x"c2"),
   465 => (x"f4",x"e0",x"c0",x"1e"),
   466 => (x"ee",x"d5",x"c2",x"1e"),
   467 => (x"87",x"cf",x"f9",x"49"),
   468 => (x"98",x"70",x"86",x"c8"),
   469 => (x"87",x"c5",x"c0",x"02"),
   470 => (x"d4",x"c3",x"48",x"c0"),
   471 => (x"dc",x"dc",x"c2",x"87"),
   472 => (x"c4",x"48",x"4a",x"bf"),
   473 => (x"ec",x"dc",x"c2",x"30"),
   474 => (x"cc",x"e1",x"c2",x"58"),
   475 => (x"c1",x"d5",x"c2",x"5a"),
   476 => (x"c8",x"49",x"bf",x"97"),
   477 => (x"c0",x"d5",x"c2",x"31"),
   478 => (x"a1",x"4b",x"bf",x"97"),
   479 => (x"c2",x"d5",x"c2",x"49"),
   480 => (x"d0",x"4b",x"bf",x"97"),
   481 => (x"49",x"a1",x"73",x"33"),
   482 => (x"97",x"c3",x"d5",x"c2"),
   483 => (x"33",x"d8",x"4b",x"bf"),
   484 => (x"c2",x"49",x"a1",x"73"),
   485 => (x"c2",x"59",x"d4",x"e1"),
   486 => (x"91",x"bf",x"cc",x"e1"),
   487 => (x"bf",x"f8",x"e0",x"c2"),
   488 => (x"c0",x"e1",x"c2",x"81"),
   489 => (x"c9",x"d5",x"c2",x"59"),
   490 => (x"c8",x"4b",x"bf",x"97"),
   491 => (x"c8",x"d5",x"c2",x"33"),
   492 => (x"a3",x"4c",x"bf",x"97"),
   493 => (x"ca",x"d5",x"c2",x"4b"),
   494 => (x"d0",x"4c",x"bf",x"97"),
   495 => (x"4b",x"a3",x"74",x"34"),
   496 => (x"97",x"cb",x"d5",x"c2"),
   497 => (x"9c",x"cf",x"4c",x"bf"),
   498 => (x"a3",x"74",x"34",x"d8"),
   499 => (x"c4",x"e1",x"c2",x"4b"),
   500 => (x"73",x"8b",x"c2",x"5b"),
   501 => (x"c4",x"e1",x"c2",x"92"),
   502 => (x"78",x"a1",x"72",x"48"),
   503 => (x"c2",x"87",x"cb",x"c1"),
   504 => (x"bf",x"97",x"ee",x"d4"),
   505 => (x"c2",x"31",x"c8",x"49"),
   506 => (x"bf",x"97",x"ed",x"d4"),
   507 => (x"c2",x"49",x"a1",x"4a"),
   508 => (x"c5",x"59",x"ec",x"dc"),
   509 => (x"81",x"ff",x"c7",x"31"),
   510 => (x"e1",x"c2",x"29",x"c9"),
   511 => (x"d4",x"c2",x"59",x"cc"),
   512 => (x"4a",x"bf",x"97",x"f3"),
   513 => (x"d4",x"c2",x"32",x"c8"),
   514 => (x"4b",x"bf",x"97",x"f2"),
   515 => (x"e1",x"c2",x"4a",x"a2"),
   516 => (x"e1",x"c2",x"5a",x"d4"),
   517 => (x"75",x"92",x"bf",x"cc"),
   518 => (x"c8",x"e1",x"c2",x"82"),
   519 => (x"c0",x"e1",x"c2",x"5a"),
   520 => (x"c2",x"78",x"c0",x"48"),
   521 => (x"72",x"48",x"fc",x"e0"),
   522 => (x"49",x"c0",x"78",x"a1"),
   523 => (x"c1",x"87",x"f7",x"c7"),
   524 => (x"87",x"e5",x"f6",x"48"),
   525 => (x"33",x"54",x"41",x"46"),
   526 => (x"20",x"20",x"20",x"32"),
   527 => (x"54",x"41",x"46",x"00"),
   528 => (x"20",x"20",x"36",x"31"),
   529 => (x"41",x"46",x"00",x"20"),
   530 => (x"20",x"32",x"33",x"54"),
   531 => (x"46",x"00",x"20",x"20"),
   532 => (x"32",x"33",x"54",x"41"),
   533 => (x"00",x"20",x"20",x"20"),
   534 => (x"31",x"54",x"41",x"46"),
   535 => (x"20",x"20",x"20",x"36"),
   536 => (x"5b",x"5e",x"0e",x"00"),
   537 => (x"71",x"0e",x"5d",x"5c"),
   538 => (x"e4",x"dc",x"c2",x"4a"),
   539 => (x"87",x"cc",x"02",x"bf"),
   540 => (x"b7",x"c7",x"4b",x"72"),
   541 => (x"c1",x"4d",x"72",x"2b"),
   542 => (x"87",x"ca",x"9d",x"ff"),
   543 => (x"b7",x"c8",x"4b",x"72"),
   544 => (x"c3",x"4d",x"72",x"2b"),
   545 => (x"d4",x"c2",x"9d",x"ff"),
   546 => (x"e0",x"c2",x"1e",x"dc"),
   547 => (x"73",x"49",x"bf",x"f8"),
   548 => (x"fe",x"ee",x"71",x"81"),
   549 => (x"70",x"86",x"c4",x"87"),
   550 => (x"87",x"c5",x"05",x"98"),
   551 => (x"e6",x"c0",x"48",x"c0"),
   552 => (x"e4",x"dc",x"c2",x"87"),
   553 => (x"87",x"d2",x"02",x"bf"),
   554 => (x"91",x"c4",x"49",x"75"),
   555 => (x"81",x"dc",x"d4",x"c2"),
   556 => (x"ff",x"cf",x"4c",x"69"),
   557 => (x"9c",x"ff",x"ff",x"ff"),
   558 => (x"49",x"75",x"87",x"cb"),
   559 => (x"d4",x"c2",x"91",x"c2"),
   560 => (x"69",x"9f",x"81",x"dc"),
   561 => (x"f4",x"48",x"74",x"4c"),
   562 => (x"5e",x"0e",x"87",x"cf"),
   563 => (x"0e",x"5d",x"5c",x"5b"),
   564 => (x"4c",x"71",x"86",x"f4"),
   565 => (x"e1",x"c2",x"4b",x"c0"),
   566 => (x"c4",x"7e",x"bf",x"d4"),
   567 => (x"e1",x"c2",x"48",x"a6"),
   568 => (x"c8",x"78",x"bf",x"d8"),
   569 => (x"78",x"c0",x"48",x"a6"),
   570 => (x"bf",x"e8",x"dc",x"c2"),
   571 => (x"06",x"a8",x"c0",x"48"),
   572 => (x"c8",x"87",x"dd",x"c2"),
   573 => (x"99",x"cf",x"49",x"66"),
   574 => (x"c2",x"87",x"d8",x"05"),
   575 => (x"c8",x"1e",x"dc",x"d4"),
   576 => (x"c1",x"48",x"49",x"66"),
   577 => (x"58",x"a6",x"cc",x"80"),
   578 => (x"c4",x"87",x"c8",x"ed"),
   579 => (x"dc",x"d4",x"c2",x"86"),
   580 => (x"c0",x"87",x"c3",x"4b"),
   581 => (x"6b",x"97",x"83",x"e0"),
   582 => (x"c1",x"02",x"9a",x"4a"),
   583 => (x"e5",x"c3",x"87",x"e1"),
   584 => (x"da",x"c1",x"02",x"aa"),
   585 => (x"49",x"a3",x"cb",x"87"),
   586 => (x"d8",x"49",x"69",x"97"),
   587 => (x"ce",x"c1",x"05",x"99"),
   588 => (x"c0",x"1e",x"cb",x"87"),
   589 => (x"73",x"1e",x"66",x"e0"),
   590 => (x"87",x"e3",x"f1",x"49"),
   591 => (x"98",x"70",x"86",x"c8"),
   592 => (x"87",x"fb",x"c0",x"05"),
   593 => (x"c4",x"4a",x"a3",x"dc"),
   594 => (x"79",x"6a",x"49",x"a4"),
   595 => (x"c8",x"49",x"a3",x"da"),
   596 => (x"69",x"9f",x"4d",x"a4"),
   597 => (x"dc",x"c2",x"7d",x"48"),
   598 => (x"d3",x"02",x"bf",x"e4"),
   599 => (x"49",x"a3",x"d4",x"87"),
   600 => (x"c0",x"49",x"69",x"9f"),
   601 => (x"71",x"99",x"ff",x"ff"),
   602 => (x"c4",x"30",x"d0",x"48"),
   603 => (x"87",x"c2",x"58",x"a6"),
   604 => (x"48",x"6e",x"7e",x"c0"),
   605 => (x"7d",x"70",x"80",x"6d"),
   606 => (x"48",x"c1",x"7c",x"c0"),
   607 => (x"c8",x"87",x"c5",x"c1"),
   608 => (x"80",x"c1",x"48",x"66"),
   609 => (x"c2",x"58",x"a6",x"cc"),
   610 => (x"a8",x"bf",x"e8",x"dc"),
   611 => (x"87",x"e3",x"fd",x"04"),
   612 => (x"bf",x"e4",x"dc",x"c2"),
   613 => (x"87",x"ea",x"c0",x"02"),
   614 => (x"c4",x"fb",x"49",x"6e"),
   615 => (x"58",x"a6",x"c4",x"87"),
   616 => (x"ff",x"cf",x"49",x"70"),
   617 => (x"99",x"f8",x"ff",x"ff"),
   618 => (x"87",x"d6",x"02",x"a9"),
   619 => (x"89",x"c2",x"49",x"70"),
   620 => (x"bf",x"dc",x"dc",x"c2"),
   621 => (x"fc",x"e0",x"c2",x"91"),
   622 => (x"80",x"71",x"48",x"bf"),
   623 => (x"fc",x"58",x"a6",x"c8"),
   624 => (x"48",x"c0",x"87",x"e1"),
   625 => (x"d0",x"f0",x"8e",x"f4"),
   626 => (x"1e",x"73",x"1e",x"87"),
   627 => (x"49",x"6a",x"4a",x"71"),
   628 => (x"7a",x"71",x"81",x"c1"),
   629 => (x"bf",x"e0",x"dc",x"c2"),
   630 => (x"87",x"cb",x"05",x"99"),
   631 => (x"6b",x"4b",x"a2",x"c8"),
   632 => (x"87",x"fd",x"f9",x"49"),
   633 => (x"c1",x"7b",x"49",x"70"),
   634 => (x"87",x"f1",x"ef",x"48"),
   635 => (x"71",x"1e",x"73",x"1e"),
   636 => (x"fc",x"e0",x"c2",x"4b"),
   637 => (x"a3",x"c8",x"49",x"bf"),
   638 => (x"c2",x"4a",x"6a",x"4a"),
   639 => (x"dc",x"dc",x"c2",x"8a"),
   640 => (x"a1",x"72",x"92",x"bf"),
   641 => (x"e0",x"dc",x"c2",x"49"),
   642 => (x"9a",x"6b",x"4a",x"bf"),
   643 => (x"c8",x"49",x"a1",x"72"),
   644 => (x"e8",x"71",x"1e",x"66"),
   645 => (x"86",x"c4",x"87",x"fd"),
   646 => (x"c4",x"05",x"98",x"70"),
   647 => (x"c2",x"48",x"c0",x"87"),
   648 => (x"ee",x"48",x"c1",x"87"),
   649 => (x"5e",x"0e",x"87",x"f7"),
   650 => (x"71",x"0e",x"5c",x"5b"),
   651 => (x"72",x"4b",x"c0",x"4a"),
   652 => (x"e0",x"c0",x"02",x"9a"),
   653 => (x"49",x"a2",x"da",x"87"),
   654 => (x"c2",x"4b",x"69",x"9f"),
   655 => (x"02",x"bf",x"e4",x"dc"),
   656 => (x"a2",x"d4",x"87",x"cf"),
   657 => (x"49",x"69",x"9f",x"49"),
   658 => (x"ff",x"ff",x"c0",x"4c"),
   659 => (x"c2",x"34",x"d0",x"9c"),
   660 => (x"74",x"4c",x"c0",x"87"),
   661 => (x"02",x"9b",x"73",x"b3"),
   662 => (x"c2",x"4a",x"87",x"df"),
   663 => (x"dc",x"dc",x"c2",x"8a"),
   664 => (x"c2",x"92",x"49",x"bf"),
   665 => (x"48",x"bf",x"fc",x"e0"),
   666 => (x"e1",x"c2",x"80",x"72"),
   667 => (x"48",x"71",x"58",x"dc"),
   668 => (x"dc",x"c2",x"30",x"c4"),
   669 => (x"e9",x"c0",x"58",x"ec"),
   670 => (x"c0",x"e1",x"c2",x"87"),
   671 => (x"e1",x"c2",x"4b",x"bf"),
   672 => (x"e1",x"c2",x"48",x"d8"),
   673 => (x"c2",x"78",x"bf",x"c4"),
   674 => (x"02",x"bf",x"e4",x"dc"),
   675 => (x"dc",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"dc"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"c8",x"e1"),
   679 => (x"dc",x"c2",x"31",x"c4"),
   680 => (x"e1",x"c2",x"59",x"ec"),
   681 => (x"f2",x"ec",x"5b",x"d8"),
   682 => (x"5b",x"5e",x"0e",x"87"),
   683 => (x"f4",x"0e",x"5d",x"5c"),
   684 => (x"9a",x"4a",x"71",x"86"),
   685 => (x"c2",x"87",x"de",x"02"),
   686 => (x"c0",x"48",x"d8",x"d4"),
   687 => (x"d0",x"d4",x"c2",x"78"),
   688 => (x"d8",x"e1",x"c2",x"48"),
   689 => (x"d4",x"c2",x"78",x"bf"),
   690 => (x"e1",x"c2",x"48",x"d4"),
   691 => (x"c0",x"78",x"bf",x"d4"),
   692 => (x"c0",x"48",x"ff",x"f1"),
   693 => (x"e8",x"dc",x"c2",x"78"),
   694 => (x"d4",x"c2",x"49",x"bf"),
   695 => (x"71",x"4a",x"bf",x"d8"),
   696 => (x"cb",x"c4",x"03",x"aa"),
   697 => (x"cf",x"49",x"72",x"87"),
   698 => (x"e0",x"c0",x"05",x"99"),
   699 => (x"dc",x"d4",x"c2",x"87"),
   700 => (x"d0",x"d4",x"c2",x"1e"),
   701 => (x"d4",x"c2",x"49",x"bf"),
   702 => (x"a1",x"c1",x"48",x"d0"),
   703 => (x"d2",x"e5",x"71",x"78"),
   704 => (x"c0",x"86",x"c4",x"87"),
   705 => (x"c2",x"48",x"fb",x"f1"),
   706 => (x"cc",x"78",x"dc",x"d4"),
   707 => (x"fb",x"f1",x"c0",x"87"),
   708 => (x"e0",x"c0",x"48",x"bf"),
   709 => (x"ff",x"f1",x"c0",x"80"),
   710 => (x"d8",x"d4",x"c2",x"58"),
   711 => (x"80",x"c1",x"48",x"bf"),
   712 => (x"58",x"dc",x"d4",x"c2"),
   713 => (x"00",x"0c",x"7b",x"27"),
   714 => (x"bf",x"97",x"bf",x"00"),
   715 => (x"c2",x"02",x"9c",x"4c"),
   716 => (x"e5",x"c3",x"87",x"ee"),
   717 => (x"e7",x"c2",x"02",x"ac"),
   718 => (x"fb",x"f1",x"c0",x"87"),
   719 => (x"a3",x"cb",x"4b",x"bf"),
   720 => (x"cf",x"4d",x"11",x"49"),
   721 => (x"d6",x"c1",x"05",x"ad"),
   722 => (x"df",x"49",x"74",x"87"),
   723 => (x"cd",x"89",x"c1",x"99"),
   724 => (x"ec",x"dc",x"c2",x"91"),
   725 => (x"4a",x"a3",x"c1",x"81"),
   726 => (x"a3",x"c3",x"51",x"12"),
   727 => (x"c5",x"51",x"12",x"4a"),
   728 => (x"51",x"12",x"4a",x"a3"),
   729 => (x"12",x"4a",x"a3",x"c7"),
   730 => (x"4a",x"a3",x"c9",x"51"),
   731 => (x"a3",x"ce",x"51",x"12"),
   732 => (x"d0",x"51",x"12",x"4a"),
   733 => (x"51",x"12",x"4a",x"a3"),
   734 => (x"12",x"4a",x"a3",x"d2"),
   735 => (x"4a",x"a3",x"d4",x"51"),
   736 => (x"a3",x"d6",x"51",x"12"),
   737 => (x"d8",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"dc"),
   740 => (x"4a",x"a3",x"de",x"51"),
   741 => (x"f1",x"c0",x"51",x"12"),
   742 => (x"78",x"c1",x"48",x"ff"),
   743 => (x"75",x"87",x"c1",x"c1"),
   744 => (x"05",x"99",x"c8",x"49"),
   745 => (x"75",x"87",x"f3",x"c0"),
   746 => (x"05",x"99",x"d0",x"49"),
   747 => (x"66",x"dc",x"87",x"d0"),
   748 => (x"87",x"ca",x"c0",x"02"),
   749 => (x"66",x"dc",x"49",x"73"),
   750 => (x"02",x"98",x"70",x"0f"),
   751 => (x"f1",x"c0",x"87",x"dc"),
   752 => (x"c0",x"05",x"bf",x"ff"),
   753 => (x"dc",x"c2",x"87",x"c6"),
   754 => (x"50",x"c0",x"48",x"ec"),
   755 => (x"48",x"ff",x"f1",x"c0"),
   756 => (x"f1",x"c0",x"78",x"c0"),
   757 => (x"c2",x"48",x"bf",x"fb"),
   758 => (x"f1",x"c0",x"87",x"dc"),
   759 => (x"78",x"c0",x"48",x"ff"),
   760 => (x"bf",x"e8",x"dc",x"c2"),
   761 => (x"d8",x"d4",x"c2",x"49"),
   762 => (x"aa",x"71",x"4a",x"bf"),
   763 => (x"87",x"f5",x"fb",x"04"),
   764 => (x"bf",x"d8",x"e1",x"c2"),
   765 => (x"87",x"c8",x"c0",x"05"),
   766 => (x"bf",x"e4",x"dc",x"c2"),
   767 => (x"87",x"f4",x"c1",x"02"),
   768 => (x"bf",x"d4",x"d4",x"c2"),
   769 => (x"87",x"d9",x"f1",x"49"),
   770 => (x"58",x"d8",x"d4",x"c2"),
   771 => (x"dc",x"c2",x"7e",x"70"),
   772 => (x"c0",x"02",x"bf",x"e4"),
   773 => (x"49",x"6e",x"87",x"dd"),
   774 => (x"ff",x"ff",x"ff",x"cf"),
   775 => (x"02",x"a9",x"99",x"f8"),
   776 => (x"c4",x"87",x"c8",x"c0"),
   777 => (x"78",x"c0",x"48",x"a6"),
   778 => (x"c4",x"87",x"e6",x"c0"),
   779 => (x"78",x"c1",x"48",x"a6"),
   780 => (x"6e",x"87",x"de",x"c0"),
   781 => (x"f8",x"ff",x"cf",x"49"),
   782 => (x"c0",x"02",x"a9",x"99"),
   783 => (x"a6",x"c8",x"87",x"c8"),
   784 => (x"c0",x"78",x"c0",x"48"),
   785 => (x"a6",x"c8",x"87",x"c5"),
   786 => (x"c4",x"78",x"c1",x"48"),
   787 => (x"66",x"c8",x"48",x"a6"),
   788 => (x"05",x"66",x"c4",x"78"),
   789 => (x"6e",x"87",x"dd",x"c0"),
   790 => (x"c2",x"89",x"c2",x"49"),
   791 => (x"91",x"bf",x"dc",x"dc"),
   792 => (x"bf",x"fc",x"e0",x"c2"),
   793 => (x"c2",x"80",x"71",x"48"),
   794 => (x"c2",x"58",x"d4",x"d4"),
   795 => (x"c0",x"48",x"d8",x"d4"),
   796 => (x"87",x"e1",x"f9",x"78"),
   797 => (x"8e",x"f4",x"48",x"c0"),
   798 => (x"00",x"87",x"de",x"e5"),
   799 => (x"00",x"00",x"00",x"00"),
   800 => (x"1e",x"00",x"00",x"00"),
   801 => (x"c3",x"48",x"d4",x"ff"),
   802 => (x"49",x"68",x"78",x"ff"),
   803 => (x"87",x"c6",x"02",x"99"),
   804 => (x"05",x"a9",x"fb",x"c0"),
   805 => (x"48",x"71",x"87",x"ee"),
   806 => (x"5e",x"0e",x"4f",x"26"),
   807 => (x"71",x"0e",x"5c",x"5b"),
   808 => (x"ff",x"4b",x"c0",x"4a"),
   809 => (x"ff",x"c3",x"48",x"d4"),
   810 => (x"99",x"49",x"68",x"78"),
   811 => (x"87",x"c1",x"c1",x"02"),
   812 => (x"02",x"a9",x"ec",x"c0"),
   813 => (x"c0",x"87",x"fa",x"c0"),
   814 => (x"c0",x"02",x"a9",x"fb"),
   815 => (x"66",x"cc",x"87",x"f3"),
   816 => (x"cc",x"03",x"ab",x"b7"),
   817 => (x"02",x"66",x"d0",x"87"),
   818 => (x"09",x"72",x"87",x"c7"),
   819 => (x"c1",x"09",x"79",x"97"),
   820 => (x"02",x"99",x"71",x"82"),
   821 => (x"83",x"c1",x"87",x"c2"),
   822 => (x"c3",x"48",x"d4",x"ff"),
   823 => (x"49",x"68",x"78",x"ff"),
   824 => (x"87",x"cd",x"02",x"99"),
   825 => (x"02",x"a9",x"ec",x"c0"),
   826 => (x"fb",x"c0",x"87",x"c7"),
   827 => (x"cd",x"ff",x"05",x"a9"),
   828 => (x"02",x"66",x"d0",x"87"),
   829 => (x"97",x"c0",x"87",x"c3"),
   830 => (x"a9",x"fb",x"c0",x"7a"),
   831 => (x"73",x"87",x"c7",x"05"),
   832 => (x"8c",x"0c",x"c0",x"4c"),
   833 => (x"4c",x"73",x"87",x"c2"),
   834 => (x"87",x"c2",x"48",x"74"),
   835 => (x"4c",x"26",x"4d",x"26"),
   836 => (x"4f",x"26",x"4b",x"26"),
   837 => (x"48",x"d4",x"ff",x"1e"),
   838 => (x"68",x"78",x"ff",x"c3"),
   839 => (x"b7",x"f0",x"c0",x"49"),
   840 => (x"87",x"ca",x"04",x"a9"),
   841 => (x"a9",x"b7",x"f9",x"c0"),
   842 => (x"c0",x"87",x"c3",x"01"),
   843 => (x"c1",x"c1",x"89",x"f0"),
   844 => (x"ca",x"04",x"a9",x"b7"),
   845 => (x"b7",x"c6",x"c1",x"87"),
   846 => (x"87",x"c3",x"01",x"a9"),
   847 => (x"71",x"89",x"f7",x"c0"),
   848 => (x"0e",x"4f",x"26",x"48"),
   849 => (x"5d",x"5c",x"5b",x"5e"),
   850 => (x"71",x"86",x"f4",x"0e"),
   851 => (x"4b",x"d4",x"ff",x"4c"),
   852 => (x"c3",x"7e",x"4d",x"c0"),
   853 => (x"d0",x"ff",x"7b",x"ff"),
   854 => (x"c0",x"c8",x"48",x"bf"),
   855 => (x"a6",x"c8",x"98",x"c0"),
   856 => (x"02",x"98",x"70",x"58"),
   857 => (x"d0",x"ff",x"87",x"d0"),
   858 => (x"c0",x"c8",x"48",x"bf"),
   859 => (x"a6",x"c8",x"98",x"c0"),
   860 => (x"05",x"98",x"70",x"58"),
   861 => (x"d0",x"ff",x"87",x"f0"),
   862 => (x"78",x"e1",x"c0",x"48"),
   863 => (x"c2",x"fc",x"7b",x"d4"),
   864 => (x"99",x"49",x"70",x"87"),
   865 => (x"87",x"c7",x"c1",x"02"),
   866 => (x"c8",x"7b",x"ff",x"c3"),
   867 => (x"78",x"6b",x"48",x"a6"),
   868 => (x"c0",x"48",x"66",x"c8"),
   869 => (x"c8",x"02",x"a8",x"fb"),
   870 => (x"f4",x"e1",x"c2",x"87"),
   871 => (x"ee",x"c0",x"02",x"bf"),
   872 => (x"71",x"4d",x"c1",x"87"),
   873 => (x"e6",x"c0",x"02",x"99"),
   874 => (x"a9",x"fb",x"c0",x"87"),
   875 => (x"fb",x"87",x"c3",x"02"),
   876 => (x"ff",x"c3",x"87",x"d1"),
   877 => (x"c1",x"49",x"6b",x"7b"),
   878 => (x"cc",x"05",x"a9",x"c6"),
   879 => (x"7b",x"ff",x"c3",x"87"),
   880 => (x"48",x"a6",x"c8",x"7b"),
   881 => (x"49",x"c0",x"78",x"6b"),
   882 => (x"05",x"99",x"71",x"4d"),
   883 => (x"75",x"87",x"da",x"ff"),
   884 => (x"de",x"c1",x"05",x"9d"),
   885 => (x"7b",x"ff",x"c3",x"87"),
   886 => (x"ff",x"c3",x"4a",x"6b"),
   887 => (x"48",x"a6",x"c4",x"7b"),
   888 => (x"48",x"6e",x"78",x"6b"),
   889 => (x"a6",x"c4",x"80",x"c1"),
   890 => (x"49",x"a4",x"c8",x"58"),
   891 => (x"c8",x"49",x"69",x"97"),
   892 => (x"da",x"05",x"a9",x"66"),
   893 => (x"49",x"a4",x"c9",x"87"),
   894 => (x"aa",x"49",x"69",x"97"),
   895 => (x"ca",x"87",x"d0",x"05"),
   896 => (x"69",x"97",x"49",x"a4"),
   897 => (x"a9",x"66",x"c4",x"49"),
   898 => (x"c1",x"87",x"c4",x"05"),
   899 => (x"c8",x"87",x"d6",x"4d"),
   900 => (x"ec",x"c0",x"48",x"66"),
   901 => (x"87",x"c9",x"02",x"a8"),
   902 => (x"c0",x"48",x"66",x"c8"),
   903 => (x"c4",x"05",x"a8",x"fb"),
   904 => (x"c1",x"7e",x"c0",x"87"),
   905 => (x"7b",x"ff",x"c3",x"4d"),
   906 => (x"6b",x"48",x"a6",x"c8"),
   907 => (x"02",x"9d",x"75",x"78"),
   908 => (x"ff",x"87",x"e2",x"fe"),
   909 => (x"c8",x"48",x"bf",x"d0"),
   910 => (x"c8",x"98",x"c0",x"c0"),
   911 => (x"98",x"70",x"58",x"a6"),
   912 => (x"ff",x"87",x"d0",x"02"),
   913 => (x"c8",x"48",x"bf",x"d0"),
   914 => (x"c8",x"98",x"c0",x"c0"),
   915 => (x"98",x"70",x"58",x"a6"),
   916 => (x"ff",x"87",x"f0",x"05"),
   917 => (x"e0",x"c0",x"48",x"d0"),
   918 => (x"f4",x"48",x"6e",x"78"),
   919 => (x"87",x"ec",x"fa",x"8e"),
   920 => (x"5c",x"5b",x"5e",x"0e"),
   921 => (x"86",x"f4",x"0e",x"5d"),
   922 => (x"ff",x"59",x"a6",x"c4"),
   923 => (x"c0",x"c8",x"4c",x"d0"),
   924 => (x"1e",x"6e",x"4b",x"c0"),
   925 => (x"49",x"f8",x"e1",x"c2"),
   926 => (x"c4",x"87",x"cf",x"e9"),
   927 => (x"02",x"98",x"70",x"86"),
   928 => (x"c2",x"87",x"f7",x"c5"),
   929 => (x"4d",x"bf",x"fc",x"e1"),
   930 => (x"f6",x"fa",x"49",x"6e"),
   931 => (x"58",x"a6",x"c8",x"87"),
   932 => (x"98",x"73",x"48",x"6c"),
   933 => (x"70",x"58",x"a6",x"cc"),
   934 => (x"87",x"cc",x"02",x"98"),
   935 => (x"98",x"73",x"48",x"6c"),
   936 => (x"70",x"58",x"a6",x"c4"),
   937 => (x"87",x"f4",x"05",x"98"),
   938 => (x"d4",x"ff",x"7c",x"c5"),
   939 => (x"78",x"d5",x"c1",x"48"),
   940 => (x"bf",x"f4",x"e1",x"c2"),
   941 => (x"c4",x"81",x"c1",x"49"),
   942 => (x"8a",x"c1",x"4a",x"66"),
   943 => (x"48",x"72",x"32",x"c6"),
   944 => (x"d4",x"ff",x"b0",x"71"),
   945 => (x"48",x"6c",x"78",x"08"),
   946 => (x"a6",x"c4",x"98",x"73"),
   947 => (x"02",x"98",x"70",x"58"),
   948 => (x"48",x"6c",x"87",x"cc"),
   949 => (x"a6",x"c4",x"98",x"73"),
   950 => (x"05",x"98",x"70",x"58"),
   951 => (x"7c",x"c4",x"87",x"f4"),
   952 => (x"c3",x"48",x"d4",x"ff"),
   953 => (x"48",x"6c",x"78",x"ff"),
   954 => (x"a6",x"c4",x"98",x"73"),
   955 => (x"02",x"98",x"70",x"58"),
   956 => (x"48",x"6c",x"87",x"cc"),
   957 => (x"a6",x"c4",x"98",x"73"),
   958 => (x"05",x"98",x"70",x"58"),
   959 => (x"7c",x"c5",x"87",x"f4"),
   960 => (x"c1",x"48",x"d4",x"ff"),
   961 => (x"78",x"c1",x"78",x"d3"),
   962 => (x"98",x"73",x"48",x"6c"),
   963 => (x"70",x"58",x"a6",x"c4"),
   964 => (x"87",x"cc",x"02",x"98"),
   965 => (x"98",x"73",x"48",x"6c"),
   966 => (x"70",x"58",x"a6",x"c4"),
   967 => (x"87",x"f4",x"05",x"98"),
   968 => (x"9d",x"75",x"7c",x"c4"),
   969 => (x"87",x"d0",x"c2",x"02"),
   970 => (x"7e",x"dc",x"d4",x"c2"),
   971 => (x"f8",x"e1",x"c2",x"1e"),
   972 => (x"87",x"f8",x"ea",x"49"),
   973 => (x"98",x"70",x"86",x"c4"),
   974 => (x"c0",x"87",x"c5",x"05"),
   975 => (x"87",x"fc",x"c2",x"48"),
   976 => (x"ad",x"b7",x"c0",x"c8"),
   977 => (x"4a",x"87",x"c4",x"04"),
   978 => (x"75",x"87",x"c4",x"8d"),
   979 => (x"6c",x"4d",x"c0",x"4a"),
   980 => (x"c8",x"98",x"73",x"48"),
   981 => (x"98",x"70",x"58",x"a6"),
   982 => (x"6c",x"87",x"cc",x"02"),
   983 => (x"c8",x"98",x"73",x"48"),
   984 => (x"98",x"70",x"58",x"a6"),
   985 => (x"cd",x"87",x"f4",x"05"),
   986 => (x"48",x"d4",x"ff",x"7c"),
   987 => (x"72",x"78",x"d4",x"c1"),
   988 => (x"71",x"8a",x"c1",x"49"),
   989 => (x"87",x"d9",x"02",x"99"),
   990 => (x"48",x"bf",x"97",x"6e"),
   991 => (x"78",x"08",x"d4",x"ff"),
   992 => (x"80",x"c1",x"48",x"6e"),
   993 => (x"72",x"58",x"a6",x"c4"),
   994 => (x"71",x"8a",x"c1",x"49"),
   995 => (x"e7",x"ff",x"05",x"99"),
   996 => (x"73",x"48",x"6c",x"87"),
   997 => (x"58",x"a6",x"c4",x"98"),
   998 => (x"cc",x"02",x"98",x"70"),
   999 => (x"73",x"48",x"6c",x"87"),
  1000 => (x"58",x"a6",x"c4",x"98"),
  1001 => (x"f4",x"05",x"98",x"70"),
  1002 => (x"c2",x"7c",x"c4",x"87"),
  1003 => (x"e8",x"49",x"f8",x"e1"),
  1004 => (x"9d",x"75",x"87",x"d7"),
  1005 => (x"87",x"f0",x"fd",x"05"),
  1006 => (x"98",x"73",x"48",x"6c"),
  1007 => (x"70",x"58",x"a6",x"c4"),
  1008 => (x"87",x"cd",x"02",x"98"),
  1009 => (x"98",x"73",x"48",x"6c"),
  1010 => (x"70",x"58",x"a6",x"c4"),
  1011 => (x"f3",x"ff",x"05",x"98"),
  1012 => (x"ff",x"7c",x"c5",x"87"),
  1013 => (x"d3",x"c1",x"48",x"d4"),
  1014 => (x"6c",x"78",x"c0",x"78"),
  1015 => (x"c4",x"98",x"73",x"48"),
  1016 => (x"98",x"70",x"58",x"a6"),
  1017 => (x"6c",x"87",x"cd",x"02"),
  1018 => (x"c4",x"98",x"73",x"48"),
  1019 => (x"98",x"70",x"58",x"a6"),
  1020 => (x"87",x"f3",x"ff",x"05"),
  1021 => (x"48",x"c1",x"7c",x"c4"),
  1022 => (x"48",x"c0",x"87",x"c2"),
  1023 => (x"cb",x"f4",x"8e",x"f4"),
  1024 => (x"5b",x"5e",x"0e",x"87"),
  1025 => (x"1e",x"0e",x"5d",x"5c"),
  1026 => (x"4c",x"c0",x"4b",x"71"),
  1027 => (x"04",x"ab",x"b7",x"4d"),
  1028 => (x"c0",x"87",x"e9",x"c0"),
  1029 => (x"75",x"1e",x"c3",x"f5"),
  1030 => (x"87",x"c4",x"02",x"9d"),
  1031 => (x"87",x"c2",x"4a",x"c0"),
  1032 => (x"49",x"72",x"4a",x"c1"),
  1033 => (x"c4",x"87",x"c2",x"ea"),
  1034 => (x"c1",x"58",x"a6",x"86"),
  1035 => (x"c2",x"05",x"6e",x"84"),
  1036 => (x"c1",x"4c",x"73",x"87"),
  1037 => (x"ac",x"b7",x"73",x"85"),
  1038 => (x"87",x"d7",x"ff",x"06"),
  1039 => (x"f3",x"26",x"48",x"6e"),
  1040 => (x"5e",x"0e",x"87",x"ca"),
  1041 => (x"0e",x"5d",x"5c",x"5b"),
  1042 => (x"c2",x"49",x"4c",x"71"),
  1043 => (x"81",x"bf",x"cc",x"e2"),
  1044 => (x"70",x"87",x"ee",x"fe"),
  1045 => (x"c0",x"02",x"9d",x"4d"),
  1046 => (x"dc",x"c2",x"87",x"f3"),
  1047 => (x"4a",x"75",x"4b",x"ec"),
  1048 => (x"c1",x"ff",x"49",x"cb"),
  1049 => (x"4b",x"74",x"87",x"ca"),
  1050 => (x"e4",x"c1",x"93",x"cb"),
  1051 => (x"83",x"c4",x"83",x"db"),
  1052 => (x"7b",x"da",x"c2",x"c1"),
  1053 => (x"c5",x"c1",x"49",x"74"),
  1054 => (x"49",x"74",x"87",x"f6"),
  1055 => (x"e2",x"c2",x"91",x"de"),
  1056 => (x"80",x"71",x"48",x"e0"),
  1057 => (x"dc",x"c2",x"7b",x"70"),
  1058 => (x"d3",x"f7",x"49",x"ec"),
  1059 => (x"c1",x"49",x"74",x"87"),
  1060 => (x"c1",x"87",x"dd",x"c5"),
  1061 => (x"f1",x"87",x"fe",x"c6"),
  1062 => (x"6f",x"4c",x"87",x"f2"),
  1063 => (x"6e",x"69",x"64",x"61"),
  1064 => (x"2e",x"2e",x"2e",x"67"),
  1065 => (x"42",x"20",x"80",x"00"),
  1066 => (x"00",x"6b",x"63",x"61"),
  1067 => (x"64",x"61",x"6f",x"4c"),
  1068 => (x"20",x"2e",x"2a",x"20"),
  1069 => (x"00",x"20",x"3a",x"00"),
  1070 => (x"61",x"42",x"20",x"80"),
  1071 => (x"80",x"00",x"6b",x"63"),
  1072 => (x"69",x"78",x"45",x"20"),
  1073 => (x"44",x"53",x"00",x"74"),
  1074 => (x"69",x"6e",x"49",x"20"),
  1075 => (x"00",x"2e",x"2e",x"74"),
  1076 => (x"42",x"00",x"4b",x"4f"),
  1077 => (x"20",x"54",x"4f",x"4f"),
  1078 => (x"52",x"20",x"20",x"20"),
  1079 => (x"1e",x"00",x"4d",x"4f"),
  1080 => (x"4b",x"71",x"1e",x"73"),
  1081 => (x"cc",x"e2",x"c2",x"49"),
  1082 => (x"d4",x"fc",x"81",x"bf"),
  1083 => (x"9a",x"4a",x"70",x"87"),
  1084 => (x"49",x"87",x"c4",x"02"),
  1085 => (x"c2",x"87",x"ef",x"e4"),
  1086 => (x"c0",x"48",x"cc",x"e2"),
  1087 => (x"c1",x"49",x"73",x"78"),
  1088 => (x"cb",x"f0",x"87",x"f8"),
  1089 => (x"1e",x"73",x"1e",x"87"),
  1090 => (x"a3",x"c4",x"4b",x"71"),
  1091 => (x"d0",x"c1",x"02",x"4a"),
  1092 => (x"02",x"8a",x"c1",x"87"),
  1093 => (x"02",x"8a",x"87",x"dc"),
  1094 => (x"8a",x"87",x"f2",x"c0"),
  1095 => (x"87",x"d3",x"c1",x"05"),
  1096 => (x"bf",x"cc",x"e2",x"c2"),
  1097 => (x"87",x"cb",x"c1",x"02"),
  1098 => (x"c2",x"88",x"c1",x"48"),
  1099 => (x"c1",x"58",x"d0",x"e2"),
  1100 => (x"e2",x"c2",x"87",x"c1"),
  1101 => (x"c6",x"49",x"bf",x"cc"),
  1102 => (x"d0",x"e2",x"c2",x"89"),
  1103 => (x"a9",x"b7",x"c0",x"59"),
  1104 => (x"87",x"ef",x"c0",x"03"),
  1105 => (x"48",x"cc",x"e2",x"c2"),
  1106 => (x"e6",x"c0",x"78",x"c0"),
  1107 => (x"c8",x"e2",x"c2",x"87"),
  1108 => (x"87",x"df",x"02",x"bf"),
  1109 => (x"bf",x"cc",x"e2",x"c2"),
  1110 => (x"c2",x"80",x"c1",x"48"),
  1111 => (x"d2",x"58",x"d0",x"e2"),
  1112 => (x"c8",x"e2",x"c2",x"87"),
  1113 => (x"87",x"cb",x"02",x"bf"),
  1114 => (x"bf",x"cc",x"e2",x"c2"),
  1115 => (x"c2",x"80",x"c6",x"48"),
  1116 => (x"73",x"58",x"d0",x"e2"),
  1117 => (x"ee",x"87",x"c3",x"49"),
  1118 => (x"5e",x"0e",x"87",x"d6"),
  1119 => (x"0e",x"5d",x"5c",x"5b"),
  1120 => (x"a6",x"d0",x"86",x"f0"),
  1121 => (x"dc",x"d4",x"c2",x"59"),
  1122 => (x"c2",x"4c",x"c0",x"4d"),
  1123 => (x"c1",x"48",x"c8",x"e2"),
  1124 => (x"48",x"a6",x"c4",x"78"),
  1125 => (x"e2",x"c2",x"78",x"c0"),
  1126 => (x"c0",x"48",x"bf",x"cc"),
  1127 => (x"c1",x"06",x"a8",x"b7"),
  1128 => (x"d4",x"c2",x"87",x"c1"),
  1129 => (x"02",x"98",x"48",x"dc"),
  1130 => (x"c0",x"87",x"f8",x"c0"),
  1131 => (x"c8",x"1e",x"c3",x"f5"),
  1132 => (x"87",x"c7",x"02",x"66"),
  1133 => (x"c0",x"48",x"a6",x"c4"),
  1134 => (x"c4",x"87",x"c5",x"78"),
  1135 => (x"78",x"c1",x"48",x"a6"),
  1136 => (x"e3",x"49",x"66",x"c4"),
  1137 => (x"86",x"c4",x"87",x"e3"),
  1138 => (x"84",x"c1",x"4d",x"70"),
  1139 => (x"c1",x"48",x"66",x"c4"),
  1140 => (x"58",x"a6",x"c8",x"80"),
  1141 => (x"bf",x"cc",x"e2",x"c2"),
  1142 => (x"c6",x"03",x"ac",x"b7"),
  1143 => (x"05",x"9d",x"75",x"87"),
  1144 => (x"c0",x"87",x"c8",x"ff"),
  1145 => (x"02",x"9d",x"75",x"4c"),
  1146 => (x"c0",x"87",x"de",x"c3"),
  1147 => (x"c8",x"1e",x"c3",x"f5"),
  1148 => (x"87",x"c7",x"02",x"66"),
  1149 => (x"c0",x"48",x"a6",x"cc"),
  1150 => (x"cc",x"87",x"c5",x"78"),
  1151 => (x"78",x"c1",x"48",x"a6"),
  1152 => (x"e2",x"49",x"66",x"cc"),
  1153 => (x"86",x"c4",x"87",x"e3"),
  1154 => (x"02",x"6e",x"58",x"a6"),
  1155 => (x"49",x"87",x"e6",x"c2"),
  1156 => (x"69",x"97",x"81",x"cb"),
  1157 => (x"02",x"99",x"d0",x"49"),
  1158 => (x"c1",x"87",x"d6",x"c1"),
  1159 => (x"74",x"4a",x"df",x"c3"),
  1160 => (x"c1",x"91",x"cb",x"49"),
  1161 => (x"72",x"81",x"db",x"e4"),
  1162 => (x"c3",x"81",x"c8",x"79"),
  1163 => (x"49",x"74",x"51",x"ff"),
  1164 => (x"e2",x"c2",x"91",x"de"),
  1165 => (x"85",x"71",x"4d",x"e0"),
  1166 => (x"7d",x"97",x"c1",x"c2"),
  1167 => (x"c0",x"49",x"a5",x"c1"),
  1168 => (x"dc",x"c2",x"51",x"e0"),
  1169 => (x"02",x"bf",x"97",x"ec"),
  1170 => (x"84",x"c1",x"87",x"d2"),
  1171 => (x"c2",x"4b",x"a5",x"c2"),
  1172 => (x"db",x"4a",x"ec",x"dc"),
  1173 => (x"d7",x"f9",x"fe",x"49"),
  1174 => (x"87",x"d9",x"c1",x"87"),
  1175 => (x"c0",x"49",x"a5",x"cd"),
  1176 => (x"c2",x"84",x"c1",x"51"),
  1177 => (x"4a",x"6e",x"4b",x"a5"),
  1178 => (x"f9",x"fe",x"49",x"cb"),
  1179 => (x"c4",x"c1",x"87",x"c2"),
  1180 => (x"cb",x"49",x"74",x"87"),
  1181 => (x"db",x"e4",x"c1",x"91"),
  1182 => (x"c2",x"c1",x"c1",x"81"),
  1183 => (x"ec",x"dc",x"c2",x"79"),
  1184 => (x"d8",x"02",x"bf",x"97"),
  1185 => (x"de",x"49",x"74",x"87"),
  1186 => (x"c2",x"84",x"c1",x"91"),
  1187 => (x"71",x"4b",x"e0",x"e2"),
  1188 => (x"ec",x"dc",x"c2",x"83"),
  1189 => (x"fe",x"49",x"dd",x"4a"),
  1190 => (x"d8",x"87",x"d5",x"f8"),
  1191 => (x"de",x"4b",x"74",x"87"),
  1192 => (x"e0",x"e2",x"c2",x"93"),
  1193 => (x"49",x"a3",x"cb",x"83"),
  1194 => (x"84",x"c1",x"51",x"c0"),
  1195 => (x"cb",x"4a",x"6e",x"73"),
  1196 => (x"fb",x"f7",x"fe",x"49"),
  1197 => (x"48",x"66",x"c4",x"87"),
  1198 => (x"a6",x"c8",x"80",x"c1"),
  1199 => (x"ac",x"b7",x"c7",x"58"),
  1200 => (x"87",x"c5",x"c0",x"03"),
  1201 => (x"e2",x"fc",x"05",x"6e"),
  1202 => (x"ac",x"b7",x"c7",x"87"),
  1203 => (x"87",x"d9",x"c0",x"03"),
  1204 => (x"48",x"c8",x"e2",x"c2"),
  1205 => (x"49",x"74",x"78",x"c0"),
  1206 => (x"e2",x"c2",x"91",x"de"),
  1207 => (x"51",x"c0",x"81",x"e0"),
  1208 => (x"b7",x"c7",x"84",x"c1"),
  1209 => (x"e7",x"ff",x"04",x"ac"),
  1210 => (x"f0",x"e5",x"c1",x"87"),
  1211 => (x"c1",x"50",x"c0",x"48"),
  1212 => (x"c1",x"48",x"e8",x"e5"),
  1213 => (x"c1",x"78",x"e1",x"cc"),
  1214 => (x"c1",x"48",x"ec",x"e5"),
  1215 => (x"c1",x"78",x"e5",x"c2"),
  1216 => (x"c1",x"48",x"f3",x"e5"),
  1217 => (x"cc",x"78",x"c5",x"c4"),
  1218 => (x"fb",x"c0",x"49",x"66"),
  1219 => (x"8e",x"f0",x"87",x"e2"),
  1220 => (x"1e",x"87",x"f9",x"e7"),
  1221 => (x"e1",x"c2",x"4a",x"71"),
  1222 => (x"49",x"72",x"5a",x"f8"),
  1223 => (x"26",x"87",x"db",x"f9"),
  1224 => (x"4a",x"71",x"1e",x"4f"),
  1225 => (x"c1",x"91",x"cb",x"49"),
  1226 => (x"c8",x"81",x"db",x"e4"),
  1227 => (x"c2",x"48",x"11",x"81"),
  1228 => (x"c0",x"58",x"f4",x"e1"),
  1229 => (x"fe",x"49",x"a2",x"f0"),
  1230 => (x"c0",x"87",x"c5",x"f6"),
  1231 => (x"87",x"d5",x"d5",x"49"),
  1232 => (x"5e",x"0e",x"4f",x"26"),
  1233 => (x"0e",x"5d",x"5c",x"5b"),
  1234 => (x"4d",x"71",x"86",x"f0"),
  1235 => (x"c1",x"91",x"cb",x"49"),
  1236 => (x"ca",x"81",x"db",x"e4"),
  1237 => (x"a6",x"c4",x"7e",x"a1"),
  1238 => (x"ec",x"e1",x"c2",x"48"),
  1239 => (x"97",x"6e",x"78",x"bf"),
  1240 => (x"66",x"c4",x"4a",x"bf"),
  1241 => (x"c8",x"2b",x"72",x"4b"),
  1242 => (x"48",x"12",x"4a",x"a1"),
  1243 => (x"70",x"58",x"a6",x"cc"),
  1244 => (x"c9",x"83",x"c1",x"9b"),
  1245 => (x"49",x"69",x"97",x"81"),
  1246 => (x"c2",x"04",x"ab",x"b7"),
  1247 => (x"6e",x"4b",x"c0",x"87"),
  1248 => (x"c8",x"4a",x"bf",x"97"),
  1249 => (x"31",x"72",x"49",x"66"),
  1250 => (x"66",x"c4",x"b9",x"ff"),
  1251 => (x"72",x"4c",x"73",x"99"),
  1252 => (x"c2",x"b4",x"71",x"34"),
  1253 => (x"ff",x"5c",x"f0",x"e1"),
  1254 => (x"ff",x"c3",x"48",x"d4"),
  1255 => (x"bf",x"d0",x"ff",x"78"),
  1256 => (x"c0",x"c0",x"c8",x"48"),
  1257 => (x"58",x"a6",x"d0",x"98"),
  1258 => (x"d0",x"02",x"98",x"70"),
  1259 => (x"bf",x"d0",x"ff",x"87"),
  1260 => (x"c0",x"c0",x"c8",x"48"),
  1261 => (x"58",x"a6",x"c4",x"98"),
  1262 => (x"f0",x"05",x"98",x"70"),
  1263 => (x"48",x"d0",x"ff",x"87"),
  1264 => (x"ff",x"78",x"e1",x"c0"),
  1265 => (x"78",x"de",x"48",x"d4"),
  1266 => (x"0c",x"7c",x"0c",x"70"),
  1267 => (x"b7",x"c8",x"48",x"74"),
  1268 => (x"08",x"d4",x"ff",x"28"),
  1269 => (x"d0",x"48",x"74",x"78"),
  1270 => (x"d4",x"ff",x"28",x"b7"),
  1271 => (x"48",x"74",x"78",x"08"),
  1272 => (x"ff",x"28",x"b7",x"d8"),
  1273 => (x"ff",x"78",x"08",x"d4"),
  1274 => (x"c8",x"48",x"bf",x"d0"),
  1275 => (x"c4",x"98",x"c0",x"c0"),
  1276 => (x"98",x"70",x"58",x"a6"),
  1277 => (x"ff",x"87",x"d0",x"02"),
  1278 => (x"c8",x"48",x"bf",x"d0"),
  1279 => (x"c4",x"98",x"c0",x"c0"),
  1280 => (x"98",x"70",x"58",x"a6"),
  1281 => (x"ff",x"87",x"f0",x"05"),
  1282 => (x"e0",x"c0",x"48",x"d0"),
  1283 => (x"c0",x"1e",x"c7",x"78"),
  1284 => (x"db",x"e4",x"c1",x"1e"),
  1285 => (x"f0",x"e1",x"c2",x"1e"),
  1286 => (x"e9",x"c1",x"49",x"bf"),
  1287 => (x"c0",x"49",x"75",x"87"),
  1288 => (x"e4",x"87",x"cd",x"f7"),
  1289 => (x"87",x"e4",x"e3",x"8e"),
  1290 => (x"71",x"1e",x"73",x"1e"),
  1291 => (x"d1",x"fc",x"49",x"4b"),
  1292 => (x"fc",x"49",x"73",x"87"),
  1293 => (x"d7",x"e3",x"87",x"cc"),
  1294 => (x"1e",x"73",x"1e",x"87"),
  1295 => (x"a3",x"c2",x"4b",x"71"),
  1296 => (x"87",x"d6",x"02",x"4a"),
  1297 => (x"c0",x"05",x"8a",x"c1"),
  1298 => (x"e2",x"c2",x"87",x"e2"),
  1299 => (x"db",x"02",x"bf",x"c4"),
  1300 => (x"88",x"c1",x"48",x"87"),
  1301 => (x"58",x"c8",x"e2",x"c2"),
  1302 => (x"e2",x"c2",x"87",x"d2"),
  1303 => (x"cb",x"02",x"bf",x"c8"),
  1304 => (x"c4",x"e2",x"c2",x"87"),
  1305 => (x"80",x"c1",x"48",x"bf"),
  1306 => (x"58",x"c8",x"e2",x"c2"),
  1307 => (x"1e",x"c0",x"1e",x"c7"),
  1308 => (x"1e",x"db",x"e4",x"c1"),
  1309 => (x"bf",x"f0",x"e1",x"c2"),
  1310 => (x"73",x"87",x"cb",x"49"),
  1311 => (x"ef",x"f5",x"c0",x"49"),
  1312 => (x"e2",x"8e",x"f4",x"87"),
  1313 => (x"5e",x"0e",x"87",x"ca"),
  1314 => (x"0e",x"5d",x"5c",x"5b"),
  1315 => (x"dc",x"86",x"d8",x"ff"),
  1316 => (x"a6",x"c8",x"59",x"a6"),
  1317 => (x"c4",x"78",x"c0",x"48"),
  1318 => (x"4d",x"78",x"c0",x"80"),
  1319 => (x"e2",x"c2",x"80",x"c4"),
  1320 => (x"c2",x"78",x"bf",x"c4"),
  1321 => (x"c1",x"48",x"c8",x"e2"),
  1322 => (x"48",x"d4",x"ff",x"78"),
  1323 => (x"ff",x"78",x"ff",x"c3"),
  1324 => (x"c8",x"48",x"bf",x"d0"),
  1325 => (x"c4",x"98",x"c0",x"c0"),
  1326 => (x"98",x"70",x"58",x"a6"),
  1327 => (x"ff",x"87",x"d0",x"02"),
  1328 => (x"c8",x"48",x"bf",x"d0"),
  1329 => (x"c4",x"98",x"c0",x"c0"),
  1330 => (x"98",x"70",x"58",x"a6"),
  1331 => (x"ff",x"87",x"f0",x"05"),
  1332 => (x"e1",x"c0",x"48",x"d0"),
  1333 => (x"48",x"d4",x"ff",x"78"),
  1334 => (x"de",x"ff",x"78",x"d4"),
  1335 => (x"d4",x"ff",x"87",x"e5"),
  1336 => (x"78",x"ff",x"c3",x"48"),
  1337 => (x"ff",x"48",x"a6",x"d4"),
  1338 => (x"d4",x"78",x"bf",x"d4"),
  1339 => (x"fb",x"c0",x"48",x"66"),
  1340 => (x"d1",x"c1",x"02",x"a8"),
  1341 => (x"66",x"f8",x"c0",x"87"),
  1342 => (x"6a",x"82",x"c4",x"4a"),
  1343 => (x"c1",x"1e",x"72",x"7e"),
  1344 => (x"c4",x"48",x"ec",x"c2"),
  1345 => (x"a1",x"c8",x"49",x"66"),
  1346 => (x"71",x"41",x"20",x"4a"),
  1347 => (x"87",x"f9",x"05",x"aa"),
  1348 => (x"4a",x"26",x"51",x"10"),
  1349 => (x"48",x"66",x"f8",x"c0"),
  1350 => (x"78",x"d3",x"cc",x"c1"),
  1351 => (x"81",x"c7",x"49",x"6a"),
  1352 => (x"c1",x"51",x"66",x"d4"),
  1353 => (x"6a",x"1e",x"d8",x"1e"),
  1354 => (x"ff",x"81",x"c8",x"49"),
  1355 => (x"c8",x"87",x"eb",x"dd"),
  1356 => (x"48",x"66",x"d0",x"86"),
  1357 => (x"01",x"a8",x"b7",x"c0"),
  1358 => (x"4d",x"c1",x"87",x"c4"),
  1359 => (x"66",x"d0",x"87",x"c8"),
  1360 => (x"d4",x"88",x"c1",x"48"),
  1361 => (x"66",x"d4",x"58",x"a6"),
  1362 => (x"87",x"e6",x"ca",x"02"),
  1363 => (x"b7",x"66",x"c0",x"c1"),
  1364 => (x"dd",x"ca",x"03",x"ad"),
  1365 => (x"48",x"d4",x"ff",x"87"),
  1366 => (x"d4",x"78",x"ff",x"c3"),
  1367 => (x"d4",x"ff",x"48",x"a6"),
  1368 => (x"66",x"d4",x"78",x"bf"),
  1369 => (x"88",x"c6",x"c1",x"48"),
  1370 => (x"70",x"58",x"a6",x"c4"),
  1371 => (x"e6",x"c0",x"02",x"98"),
  1372 => (x"88",x"c9",x"48",x"87"),
  1373 => (x"70",x"58",x"a6",x"c4"),
  1374 => (x"ce",x"c4",x"02",x"98"),
  1375 => (x"88",x"c1",x"48",x"87"),
  1376 => (x"70",x"58",x"a6",x"c4"),
  1377 => (x"e0",x"c1",x"02",x"98"),
  1378 => (x"88",x"c4",x"48",x"87"),
  1379 => (x"98",x"70",x"58",x"a6"),
  1380 => (x"87",x"f7",x"c3",x"02"),
  1381 => (x"d8",x"87",x"c5",x"c9"),
  1382 => (x"c2",x"c1",x"05",x"66"),
  1383 => (x"48",x"d4",x"ff",x"87"),
  1384 => (x"c0",x"78",x"ff",x"c3"),
  1385 => (x"75",x"1e",x"ca",x"1e"),
  1386 => (x"c1",x"93",x"cb",x"4b"),
  1387 => (x"c4",x"83",x"66",x"c0"),
  1388 => (x"49",x"6c",x"4c",x"a3"),
  1389 => (x"87",x"e2",x"db",x"ff"),
  1390 => (x"1e",x"de",x"1e",x"c1"),
  1391 => (x"db",x"ff",x"49",x"6c"),
  1392 => (x"86",x"d0",x"87",x"d8"),
  1393 => (x"7b",x"d3",x"cc",x"c1"),
  1394 => (x"ad",x"b7",x"66",x"d0"),
  1395 => (x"c1",x"87",x"c5",x"04"),
  1396 => (x"87",x"cf",x"c8",x"85"),
  1397 => (x"c1",x"48",x"66",x"d0"),
  1398 => (x"58",x"a6",x"d4",x"88"),
  1399 => (x"ff",x"87",x"c4",x"c8"),
  1400 => (x"d8",x"87",x"e0",x"da"),
  1401 => (x"fa",x"c7",x"58",x"a6"),
  1402 => (x"e7",x"dc",x"ff",x"87"),
  1403 => (x"58",x"a6",x"cc",x"87"),
  1404 => (x"a8",x"b7",x"66",x"cc"),
  1405 => (x"cc",x"87",x"c6",x"06"),
  1406 => (x"66",x"c8",x"48",x"a6"),
  1407 => (x"d3",x"dc",x"ff",x"78"),
  1408 => (x"a8",x"ec",x"c0",x"87"),
  1409 => (x"87",x"c3",x"c2",x"05"),
  1410 => (x"c1",x"05",x"66",x"d8"),
  1411 => (x"49",x"75",x"87",x"f3"),
  1412 => (x"f8",x"c0",x"91",x"cb"),
  1413 => (x"a1",x"c4",x"81",x"66"),
  1414 => (x"c8",x"4c",x"6a",x"4a"),
  1415 => (x"66",x"c8",x"4a",x"a1"),
  1416 => (x"e1",x"cc",x"c1",x"52"),
  1417 => (x"48",x"d4",x"ff",x"79"),
  1418 => (x"d4",x"78",x"ff",x"c3"),
  1419 => (x"d4",x"ff",x"48",x"a6"),
  1420 => (x"66",x"d4",x"78",x"bf"),
  1421 => (x"87",x"e8",x"c0",x"02"),
  1422 => (x"a8",x"fb",x"c0",x"48"),
  1423 => (x"87",x"e0",x"c0",x"02"),
  1424 => (x"7c",x"97",x"66",x"d4"),
  1425 => (x"d4",x"ff",x"84",x"c1"),
  1426 => (x"78",x"ff",x"c3",x"48"),
  1427 => (x"ff",x"48",x"a6",x"d4"),
  1428 => (x"d4",x"78",x"bf",x"d4"),
  1429 => (x"87",x"c8",x"02",x"66"),
  1430 => (x"a8",x"fb",x"c0",x"48"),
  1431 => (x"87",x"e0",x"ff",x"05"),
  1432 => (x"c2",x"54",x"e0",x"c0"),
  1433 => (x"97",x"c0",x"54",x"c1"),
  1434 => (x"b7",x"66",x"d0",x"7c"),
  1435 => (x"c5",x"c0",x"04",x"ad"),
  1436 => (x"c5",x"85",x"c1",x"87"),
  1437 => (x"66",x"d0",x"87",x"ed"),
  1438 => (x"d4",x"88",x"c1",x"48"),
  1439 => (x"e2",x"c5",x"58",x"a6"),
  1440 => (x"fe",x"d7",x"ff",x"87"),
  1441 => (x"58",x"a6",x"d8",x"87"),
  1442 => (x"c8",x"87",x"d8",x"c5"),
  1443 => (x"66",x"d8",x"48",x"66"),
  1444 => (x"fd",x"c4",x"05",x"a8"),
  1445 => (x"48",x"a6",x"dc",x"87"),
  1446 => (x"d9",x"ff",x"78",x"c0"),
  1447 => (x"a6",x"d8",x"87",x"f6"),
  1448 => (x"ef",x"d9",x"ff",x"58"),
  1449 => (x"a6",x"e4",x"c0",x"87"),
  1450 => (x"a8",x"ec",x"c0",x"58"),
  1451 => (x"87",x"ca",x"c0",x"05"),
  1452 => (x"48",x"a6",x"e0",x"c0"),
  1453 => (x"c0",x"78",x"66",x"d4"),
  1454 => (x"d4",x"ff",x"87",x"c6"),
  1455 => (x"78",x"ff",x"c3",x"48"),
  1456 => (x"91",x"cb",x"49",x"75"),
  1457 => (x"48",x"66",x"f8",x"c0"),
  1458 => (x"a6",x"c4",x"80",x"71"),
  1459 => (x"ca",x"49",x"6e",x"58"),
  1460 => (x"51",x"66",x"d4",x"81"),
  1461 => (x"49",x"66",x"e0",x"c0"),
  1462 => (x"66",x"d4",x"81",x"c1"),
  1463 => (x"71",x"48",x"c1",x"89"),
  1464 => (x"c1",x"49",x"70",x"30"),
  1465 => (x"c8",x"4a",x"6e",x"89"),
  1466 => (x"97",x"09",x"72",x"82"),
  1467 => (x"e1",x"c2",x"09",x"79"),
  1468 => (x"d4",x"49",x"bf",x"ec"),
  1469 => (x"97",x"29",x"b7",x"66"),
  1470 => (x"71",x"48",x"4a",x"6a"),
  1471 => (x"a6",x"e8",x"c0",x"98"),
  1472 => (x"c4",x"48",x"6e",x"58"),
  1473 => (x"58",x"a6",x"c8",x"80"),
  1474 => (x"4c",x"bf",x"66",x"c4"),
  1475 => (x"c8",x"48",x"66",x"d8"),
  1476 => (x"c0",x"02",x"a8",x"66"),
  1477 => (x"e0",x"c0",x"87",x"c9"),
  1478 => (x"78",x"c0",x"48",x"a6"),
  1479 => (x"c0",x"87",x"c6",x"c0"),
  1480 => (x"c1",x"48",x"a6",x"e0"),
  1481 => (x"66",x"e0",x"c0",x"78"),
  1482 => (x"1e",x"e0",x"c0",x"1e"),
  1483 => (x"d5",x"ff",x"49",x"74"),
  1484 => (x"86",x"c8",x"87",x"e8"),
  1485 => (x"c0",x"58",x"a6",x"d8"),
  1486 => (x"c1",x"06",x"a8",x"b7"),
  1487 => (x"66",x"d4",x"87",x"da"),
  1488 => (x"bf",x"66",x"c4",x"84"),
  1489 => (x"81",x"e0",x"c0",x"49"),
  1490 => (x"c1",x"4b",x"89",x"74"),
  1491 => (x"71",x"4a",x"f5",x"c2"),
  1492 => (x"87",x"dc",x"e5",x"fe"),
  1493 => (x"66",x"dc",x"84",x"c2"),
  1494 => (x"c0",x"80",x"c1",x"48"),
  1495 => (x"c0",x"58",x"a6",x"e0"),
  1496 => (x"c1",x"49",x"66",x"e4"),
  1497 => (x"02",x"a9",x"70",x"81"),
  1498 => (x"c0",x"87",x"c9",x"c0"),
  1499 => (x"c0",x"48",x"a6",x"e0"),
  1500 => (x"87",x"c6",x"c0",x"78"),
  1501 => (x"48",x"a6",x"e0",x"c0"),
  1502 => (x"e0",x"c0",x"78",x"c1"),
  1503 => (x"66",x"c8",x"1e",x"66"),
  1504 => (x"e0",x"c0",x"49",x"bf"),
  1505 => (x"71",x"89",x"74",x"81"),
  1506 => (x"ff",x"49",x"74",x"1e"),
  1507 => (x"c8",x"87",x"cb",x"d4"),
  1508 => (x"a8",x"b7",x"c0",x"86"),
  1509 => (x"87",x"fe",x"fe",x"01"),
  1510 => (x"c0",x"02",x"66",x"dc"),
  1511 => (x"49",x"6e",x"87",x"d0"),
  1512 => (x"66",x"dc",x"81",x"c9"),
  1513 => (x"c1",x"48",x"6e",x"51"),
  1514 => (x"c0",x"78",x"c2",x"cd"),
  1515 => (x"49",x"6e",x"87",x"cc"),
  1516 => (x"51",x"c2",x"81",x"c9"),
  1517 => (x"d0",x"c1",x"48",x"6e"),
  1518 => (x"66",x"d0",x"78",x"e8"),
  1519 => (x"c0",x"04",x"ad",x"b7"),
  1520 => (x"85",x"c1",x"87",x"c5"),
  1521 => (x"d0",x"87",x"dc",x"c0"),
  1522 => (x"88",x"c1",x"48",x"66"),
  1523 => (x"c0",x"58",x"a6",x"d4"),
  1524 => (x"d2",x"ff",x"87",x"d1"),
  1525 => (x"a6",x"d8",x"87",x"ed"),
  1526 => (x"87",x"c7",x"c0",x"58"),
  1527 => (x"87",x"e3",x"d2",x"ff"),
  1528 => (x"d4",x"58",x"a6",x"d8"),
  1529 => (x"c9",x"c0",x"02",x"66"),
  1530 => (x"66",x"c0",x"c1",x"87"),
  1531 => (x"f5",x"04",x"ad",x"b7"),
  1532 => (x"b7",x"c7",x"87",x"e3"),
  1533 => (x"df",x"c0",x"03",x"ad"),
  1534 => (x"c8",x"e2",x"c2",x"87"),
  1535 => (x"75",x"78",x"c0",x"48"),
  1536 => (x"c0",x"91",x"cb",x"49"),
  1537 => (x"c4",x"81",x"66",x"f8"),
  1538 => (x"4a",x"6a",x"4a",x"a1"),
  1539 => (x"c1",x"79",x"52",x"c0"),
  1540 => (x"ad",x"b7",x"c7",x"85"),
  1541 => (x"87",x"e1",x"ff",x"04"),
  1542 => (x"c0",x"02",x"66",x"d8"),
  1543 => (x"f8",x"c0",x"87",x"e2"),
  1544 => (x"cd",x"c1",x"49",x"66"),
  1545 => (x"66",x"f8",x"c0",x"81"),
  1546 => (x"82",x"d5",x"c1",x"4a"),
  1547 => (x"cc",x"c1",x"52",x"c0"),
  1548 => (x"f8",x"c0",x"79",x"e1"),
  1549 => (x"d1",x"c1",x"49",x"66"),
  1550 => (x"f8",x"c2",x"c1",x"81"),
  1551 => (x"87",x"d6",x"c0",x"79"),
  1552 => (x"49",x"66",x"f8",x"c0"),
  1553 => (x"c0",x"81",x"cd",x"c1"),
  1554 => (x"c1",x"4a",x"66",x"f8"),
  1555 => (x"c2",x"c1",x"82",x"d1"),
  1556 => (x"c9",x"c2",x"7a",x"ff"),
  1557 => (x"d0",x"c1",x"79",x"d5"),
  1558 => (x"f8",x"c0",x"4a",x"f9"),
  1559 => (x"d8",x"c1",x"49",x"66"),
  1560 => (x"ff",x"79",x"72",x"81"),
  1561 => (x"c8",x"48",x"bf",x"d0"),
  1562 => (x"c4",x"98",x"c0",x"c0"),
  1563 => (x"98",x"70",x"58",x"a6"),
  1564 => (x"87",x"d1",x"c0",x"02"),
  1565 => (x"48",x"bf",x"d0",x"ff"),
  1566 => (x"98",x"c0",x"c0",x"c8"),
  1567 => (x"70",x"58",x"a6",x"c4"),
  1568 => (x"ef",x"ff",x"05",x"98"),
  1569 => (x"48",x"d0",x"ff",x"87"),
  1570 => (x"cc",x"78",x"e0",x"c0"),
  1571 => (x"d8",x"ff",x"48",x"66"),
  1572 => (x"f7",x"d1",x"ff",x"8e"),
  1573 => (x"1e",x"c7",x"1e",x"87"),
  1574 => (x"e4",x"c1",x"1e",x"c0"),
  1575 => (x"e1",x"c2",x"1e",x"db"),
  1576 => (x"ef",x"49",x"bf",x"f0"),
  1577 => (x"e4",x"c1",x"87",x"e0"),
  1578 => (x"e6",x"c0",x"49",x"db"),
  1579 => (x"8e",x"f4",x"87",x"d4"),
  1580 => (x"c9",x"1e",x"4f",x"26"),
  1581 => (x"e2",x"c2",x"87",x"fd"),
  1582 => (x"50",x"c0",x"48",x"d0"),
  1583 => (x"c3",x"48",x"d4",x"ff"),
  1584 => (x"c3",x"c1",x"78",x"ff"),
  1585 => (x"df",x"fe",x"49",x"c6"),
  1586 => (x"e8",x"fe",x"87",x"c2"),
  1587 => (x"98",x"70",x"87",x"cd"),
  1588 => (x"fe",x"87",x"cd",x"02"),
  1589 => (x"70",x"87",x"ca",x"f4"),
  1590 => (x"87",x"c4",x"02",x"98"),
  1591 => (x"87",x"c2",x"4a",x"c1"),
  1592 => (x"9a",x"72",x"4a",x"c0"),
  1593 => (x"c1",x"87",x"c8",x"02"),
  1594 => (x"fe",x"49",x"d0",x"c3"),
  1595 => (x"c2",x"87",x"dd",x"de"),
  1596 => (x"49",x"bf",x"dc",x"d3"),
  1597 => (x"87",x"e8",x"d5",x"ff"),
  1598 => (x"48",x"c4",x"e2",x"c2"),
  1599 => (x"e1",x"c2",x"78",x"c0"),
  1600 => (x"78",x"c0",x"48",x"f0"),
  1601 => (x"87",x"cd",x"fe",x"49"),
  1602 => (x"c8",x"87",x"d4",x"c3"),
  1603 => (x"e5",x"c0",x"87",x"f9"),
  1604 => (x"f6",x"ff",x"87",x"d2"),
  1605 => (x"d3",x"4f",x"26",x"87"),
  1606 => (x"42",x"00",x"00",x"10"),
  1607 => (x"a0",x"00",x"00",x"10"),
  1608 => (x"00",x"00",x"00",x"28"),
  1609 => (x"10",x"42",x"00",x"00"),
  1610 => (x"28",x"be",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"10",x"42",x"00"),
  1613 => (x"00",x"28",x"dc",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"10",x"42"),
  1616 => (x"00",x"00",x"28",x"fa"),
  1617 => (x"42",x"00",x"00",x"00"),
  1618 => (x"18",x"00",x"00",x"10"),
  1619 => (x"00",x"00",x"00",x"29"),
  1620 => (x"10",x"42",x"00",x"00"),
  1621 => (x"29",x"36",x"00",x"00"),
  1622 => (x"00",x"00",x"00",x"00"),
  1623 => (x"00",x"10",x"42",x"00"),
  1624 => (x"00",x"29",x"54",x"00"),
  1625 => (x"00",x"00",x"00",x"00"),
  1626 => (x"00",x"00",x"13",x"21"),
  1627 => (x"00",x"00",x"00",x"00"),
  1628 => (x"05",x"00",x"00",x"00"),
  1629 => (x"00",x"00",x"00",x"11"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"1e",x"1e",x"00",x"00"),
  1632 => (x"c4",x"87",x"d5",x"c1"),
  1633 => (x"26",x"26",x"58",x"a6"),
  1634 => (x"4a",x"71",x"1e",x"4f"),
  1635 => (x"c0",x"48",x"f0",x"fe"),
  1636 => (x"7a",x"0a",x"cd",x"78"),
  1637 => (x"df",x"e6",x"c1",x"0a"),
  1638 => (x"ef",x"db",x"fe",x"49"),
  1639 => (x"53",x"4f",x"26",x"87"),
  1640 => (x"68",x"20",x"74",x"65"),
  1641 => (x"6c",x"64",x"6e",x"61"),
  1642 => (x"00",x"0a",x"72",x"65"),
  1643 => (x"69",x"20",x"6e",x"49"),
  1644 => (x"72",x"65",x"74",x"6e"),
  1645 => (x"74",x"70",x"75",x"72"),
  1646 => (x"6e",x"6f",x"63",x"20"),
  1647 => (x"75",x"72",x"74",x"73"),
  1648 => (x"72",x"6f",x"74",x"63"),
  1649 => (x"c1",x"1e",x"00",x"0a"),
  1650 => (x"fe",x"49",x"ec",x"e6"),
  1651 => (x"c1",x"87",x"fd",x"da"),
  1652 => (x"fe",x"49",x"fe",x"e5"),
  1653 => (x"4f",x"26",x"87",x"f3"),
  1654 => (x"bf",x"f0",x"fe",x"1e"),
  1655 => (x"1e",x"4f",x"26",x"48"),
  1656 => (x"c1",x"48",x"f0",x"fe"),
  1657 => (x"1e",x"4f",x"26",x"78"),
  1658 => (x"c0",x"48",x"f0",x"fe"),
  1659 => (x"1e",x"4f",x"26",x"78"),
  1660 => (x"7a",x"c0",x"4a",x"71"),
  1661 => (x"c0",x"49",x"a2",x"c4"),
  1662 => (x"49",x"a2",x"c8",x"79"),
  1663 => (x"a2",x"cc",x"79",x"c0"),
  1664 => (x"26",x"79",x"c0",x"49"),
  1665 => (x"5b",x"5e",x"0e",x"4f"),
  1666 => (x"86",x"f8",x"0e",x"5c"),
  1667 => (x"a4",x"c8",x"4c",x"71"),
  1668 => (x"4b",x"a4",x"cc",x"49"),
  1669 => (x"80",x"c1",x"48",x"6b"),
  1670 => (x"cf",x"58",x"a6",x"c4"),
  1671 => (x"58",x"a6",x"c8",x"98"),
  1672 => (x"66",x"c4",x"48",x"69"),
  1673 => (x"87",x"d4",x"05",x"a8"),
  1674 => (x"80",x"c1",x"48",x"6b"),
  1675 => (x"cf",x"58",x"a6",x"c4"),
  1676 => (x"58",x"a6",x"c8",x"98"),
  1677 => (x"66",x"c4",x"48",x"69"),
  1678 => (x"87",x"ec",x"02",x"a8"),
  1679 => (x"c1",x"87",x"e8",x"fe"),
  1680 => (x"6b",x"49",x"a4",x"d0"),
  1681 => (x"c4",x"90",x"c4",x"48"),
  1682 => (x"81",x"70",x"58",x"a6"),
  1683 => (x"6b",x"79",x"66",x"d4"),
  1684 => (x"c8",x"80",x"c1",x"48"),
  1685 => (x"98",x"cf",x"58",x"a6"),
  1686 => (x"d2",x"c1",x"7b",x"70"),
  1687 => (x"87",x"ff",x"fd",x"87"),
  1688 => (x"87",x"c2",x"8e",x"f8"),
  1689 => (x"4c",x"26",x"4d",x"26"),
  1690 => (x"4f",x"26",x"4b",x"26"),
  1691 => (x"5c",x"5b",x"5e",x"0e"),
  1692 => (x"86",x"f8",x"0e",x"5d"),
  1693 => (x"a5",x"c4",x"4d",x"71"),
  1694 => (x"6c",x"48",x"6d",x"4c"),
  1695 => (x"87",x"c5",x"05",x"a8"),
  1696 => (x"e5",x"c0",x"48",x"ff"),
  1697 => (x"87",x"df",x"fd",x"87"),
  1698 => (x"6c",x"4b",x"a5",x"d0"),
  1699 => (x"c4",x"90",x"c4",x"48"),
  1700 => (x"83",x"70",x"58",x"a6"),
  1701 => (x"ff",x"c3",x"4b",x"6b"),
  1702 => (x"c1",x"48",x"6c",x"9b"),
  1703 => (x"58",x"a6",x"c8",x"80"),
  1704 => (x"7c",x"70",x"98",x"cf"),
  1705 => (x"73",x"87",x"f8",x"fc"),
  1706 => (x"8e",x"f8",x"48",x"49"),
  1707 => (x"1e",x"87",x"f5",x"fe"),
  1708 => (x"86",x"f8",x"1e",x"73"),
  1709 => (x"e0",x"87",x"f0",x"fc"),
  1710 => (x"c0",x"49",x"4b",x"bf"),
  1711 => (x"02",x"99",x"c0",x"e0"),
  1712 => (x"73",x"87",x"e7",x"c0"),
  1713 => (x"9a",x"ff",x"c3",x"4a"),
  1714 => (x"bf",x"f2",x"e5",x"c2"),
  1715 => (x"c4",x"90",x"c4",x"48"),
  1716 => (x"e6",x"c2",x"58",x"a6"),
  1717 => (x"81",x"70",x"49",x"c2"),
  1718 => (x"e5",x"c2",x"79",x"72"),
  1719 => (x"c1",x"48",x"bf",x"f2"),
  1720 => (x"58",x"a6",x"c8",x"80"),
  1721 => (x"e5",x"c2",x"98",x"cf"),
  1722 => (x"49",x"73",x"58",x"f6"),
  1723 => (x"02",x"99",x"c0",x"d0"),
  1724 => (x"c2",x"87",x"f2",x"c0"),
  1725 => (x"48",x"bf",x"fa",x"e5"),
  1726 => (x"bf",x"fe",x"e5",x"c2"),
  1727 => (x"e4",x"c0",x"02",x"a8"),
  1728 => (x"fa",x"e5",x"c2",x"87"),
  1729 => (x"90",x"c4",x"48",x"bf"),
  1730 => (x"c2",x"58",x"a6",x"c4"),
  1731 => (x"70",x"49",x"c2",x"e7"),
  1732 => (x"69",x"48",x"e0",x"81"),
  1733 => (x"fa",x"e5",x"c2",x"78"),
  1734 => (x"80",x"c1",x"48",x"bf"),
  1735 => (x"cf",x"58",x"a6",x"c8"),
  1736 => (x"fe",x"e5",x"c2",x"98"),
  1737 => (x"87",x"f0",x"fa",x"58"),
  1738 => (x"fa",x"58",x"a6",x"c4"),
  1739 => (x"8e",x"f8",x"87",x"f1"),
  1740 => (x"1e",x"87",x"f5",x"fc"),
  1741 => (x"49",x"f2",x"e5",x"c2"),
  1742 => (x"c1",x"87",x"f4",x"fa"),
  1743 => (x"f9",x"49",x"ef",x"ea"),
  1744 => (x"f5",x"c3",x"87",x"c7"),
  1745 => (x"1e",x"4f",x"26",x"87"),
  1746 => (x"e5",x"c2",x"1e",x"73"),
  1747 => (x"db",x"fc",x"49",x"f2"),
  1748 => (x"c0",x"4a",x"70",x"87"),
  1749 => (x"c2",x"04",x"aa",x"b7"),
  1750 => (x"f0",x"c3",x"87",x"cc"),
  1751 => (x"87",x"c9",x"05",x"aa"),
  1752 => (x"48",x"f2",x"ef",x"c1"),
  1753 => (x"ed",x"c1",x"78",x"c1"),
  1754 => (x"aa",x"e0",x"c3",x"87"),
  1755 => (x"c1",x"87",x"c9",x"05"),
  1756 => (x"c1",x"48",x"f6",x"ef"),
  1757 => (x"87",x"de",x"c1",x"78"),
  1758 => (x"bf",x"f6",x"ef",x"c1"),
  1759 => (x"c2",x"87",x"c6",x"02"),
  1760 => (x"c2",x"4b",x"a2",x"c0"),
  1761 => (x"c1",x"4b",x"72",x"87"),
  1762 => (x"02",x"bf",x"f2",x"ef"),
  1763 => (x"73",x"87",x"e0",x"c0"),
  1764 => (x"29",x"b7",x"c4",x"49"),
  1765 => (x"fa",x"ef",x"c1",x"91"),
  1766 => (x"cf",x"4a",x"73",x"81"),
  1767 => (x"c1",x"92",x"c2",x"9a"),
  1768 => (x"70",x"30",x"72",x"48"),
  1769 => (x"72",x"ba",x"ff",x"4a"),
  1770 => (x"70",x"98",x"69",x"48"),
  1771 => (x"73",x"87",x"db",x"79"),
  1772 => (x"29",x"b7",x"c4",x"49"),
  1773 => (x"fa",x"ef",x"c1",x"91"),
  1774 => (x"cf",x"4a",x"73",x"81"),
  1775 => (x"c3",x"92",x"c2",x"9a"),
  1776 => (x"70",x"30",x"72",x"48"),
  1777 => (x"b0",x"69",x"48",x"4a"),
  1778 => (x"ef",x"c1",x"79",x"70"),
  1779 => (x"78",x"c0",x"48",x"f6"),
  1780 => (x"48",x"f2",x"ef",x"c1"),
  1781 => (x"e5",x"c2",x"78",x"c0"),
  1782 => (x"cf",x"fa",x"49",x"f2"),
  1783 => (x"c0",x"4a",x"70",x"87"),
  1784 => (x"fd",x"03",x"aa",x"b7"),
  1785 => (x"48",x"c0",x"87",x"f4"),
  1786 => (x"4d",x"26",x"87",x"c4"),
  1787 => (x"4b",x"26",x"4c",x"26"),
  1788 => (x"00",x"00",x"4f",x"26"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"c0",x"1e",x"00",x"00"),
  1807 => (x"c4",x"49",x"72",x"4a"),
  1808 => (x"fa",x"ef",x"c1",x"91"),
  1809 => (x"c1",x"79",x"c0",x"81"),
  1810 => (x"aa",x"b7",x"d0",x"82"),
  1811 => (x"26",x"87",x"ee",x"04"),
  1812 => (x"5b",x"5e",x"0e",x"4f"),
  1813 => (x"71",x"0e",x"5d",x"5c"),
  1814 => (x"87",x"cb",x"f6",x"4d"),
  1815 => (x"b7",x"c4",x"4a",x"75"),
  1816 => (x"ef",x"c1",x"92",x"2a"),
  1817 => (x"4c",x"75",x"82",x"fa"),
  1818 => (x"94",x"c2",x"9c",x"cf"),
  1819 => (x"74",x"4b",x"49",x"6a"),
  1820 => (x"c2",x"9b",x"c3",x"2b"),
  1821 => (x"70",x"30",x"74",x"48"),
  1822 => (x"74",x"bc",x"ff",x"4c"),
  1823 => (x"70",x"98",x"71",x"48"),
  1824 => (x"87",x"db",x"f5",x"7a"),
  1825 => (x"e1",x"fd",x"48",x"73"),
  1826 => (x"ff",x"1e",x"1e",x"87"),
  1827 => (x"c8",x"48",x"bf",x"d0"),
  1828 => (x"c4",x"98",x"c0",x"c0"),
  1829 => (x"98",x"70",x"58",x"a6"),
  1830 => (x"ff",x"87",x"d0",x"02"),
  1831 => (x"c8",x"48",x"bf",x"d0"),
  1832 => (x"c4",x"98",x"c0",x"c0"),
  1833 => (x"98",x"70",x"58",x"a6"),
  1834 => (x"ff",x"87",x"f0",x"05"),
  1835 => (x"e1",x"c4",x"48",x"d0"),
  1836 => (x"ff",x"48",x"71",x"78"),
  1837 => (x"c8",x"78",x"08",x"d4"),
  1838 => (x"d4",x"ff",x"48",x"66"),
  1839 => (x"26",x"26",x"78",x"08"),
  1840 => (x"71",x"1e",x"1e",x"4f"),
  1841 => (x"49",x"66",x"c8",x"4a"),
  1842 => (x"fe",x"49",x"72",x"1e"),
  1843 => (x"86",x"c4",x"87",x"fb"),
  1844 => (x"48",x"bf",x"d0",x"ff"),
  1845 => (x"98",x"c0",x"c0",x"c8"),
  1846 => (x"70",x"58",x"a6",x"c4"),
  1847 => (x"87",x"d0",x"02",x"98"),
  1848 => (x"48",x"bf",x"d0",x"ff"),
  1849 => (x"98",x"c0",x"c0",x"c8"),
  1850 => (x"70",x"58",x"a6",x"c4"),
  1851 => (x"87",x"f0",x"05",x"98"),
  1852 => (x"c0",x"48",x"d0",x"ff"),
  1853 => (x"26",x"26",x"78",x"e0"),
  1854 => (x"1e",x"73",x"1e",x"4f"),
  1855 => (x"66",x"c8",x"4b",x"71"),
  1856 => (x"c1",x"4a",x"73",x"1e"),
  1857 => (x"fe",x"49",x"a2",x"e0"),
  1858 => (x"c4",x"26",x"87",x"f7"),
  1859 => (x"26",x"4d",x"26",x"87"),
  1860 => (x"26",x"4b",x"26",x"4c"),
  1861 => (x"ff",x"1e",x"1e",x"4f"),
  1862 => (x"c8",x"48",x"bf",x"d0"),
  1863 => (x"c4",x"98",x"c0",x"c0"),
  1864 => (x"98",x"70",x"58",x"a6"),
  1865 => (x"ff",x"87",x"d0",x"02"),
  1866 => (x"c8",x"48",x"bf",x"d0"),
  1867 => (x"c4",x"98",x"c0",x"c0"),
  1868 => (x"98",x"70",x"58",x"a6"),
  1869 => (x"ff",x"87",x"f0",x"05"),
  1870 => (x"c9",x"c4",x"48",x"d0"),
  1871 => (x"ff",x"48",x"71",x"78"),
  1872 => (x"26",x"78",x"08",x"d4"),
  1873 => (x"1e",x"1e",x"4f",x"26"),
  1874 => (x"ff",x"49",x"4a",x"71"),
  1875 => (x"d0",x"ff",x"87",x"c7"),
  1876 => (x"c0",x"c8",x"48",x"bf"),
  1877 => (x"a6",x"c4",x"98",x"c0"),
  1878 => (x"02",x"98",x"70",x"58"),
  1879 => (x"d0",x"ff",x"87",x"d0"),
  1880 => (x"c0",x"c8",x"48",x"bf"),
  1881 => (x"a6",x"c4",x"98",x"c0"),
  1882 => (x"05",x"98",x"70",x"58"),
  1883 => (x"d0",x"ff",x"87",x"f0"),
  1884 => (x"26",x"78",x"c8",x"48"),
  1885 => (x"73",x"1e",x"4f",x"26"),
  1886 => (x"4b",x"71",x"1e",x"1e"),
  1887 => (x"bf",x"ce",x"e8",x"c2"),
  1888 => (x"c3",x"87",x"c3",x"02"),
  1889 => (x"d0",x"ff",x"87",x"cc"),
  1890 => (x"c0",x"c8",x"48",x"bf"),
  1891 => (x"a6",x"c4",x"98",x"c0"),
  1892 => (x"02",x"98",x"70",x"58"),
  1893 => (x"d0",x"ff",x"87",x"d0"),
  1894 => (x"c0",x"c8",x"48",x"bf"),
  1895 => (x"a6",x"c4",x"98",x"c0"),
  1896 => (x"05",x"98",x"70",x"58"),
  1897 => (x"d0",x"ff",x"87",x"f0"),
  1898 => (x"78",x"c9",x"c4",x"48"),
  1899 => (x"e0",x"c0",x"48",x"73"),
  1900 => (x"08",x"d4",x"ff",x"b0"),
  1901 => (x"c2",x"e8",x"c2",x"78"),
  1902 => (x"cc",x"78",x"c0",x"48"),
  1903 => (x"87",x"c5",x"02",x"66"),
  1904 => (x"c2",x"49",x"ff",x"c3"),
  1905 => (x"c2",x"49",x"c0",x"87"),
  1906 => (x"d0",x"59",x"ca",x"e8"),
  1907 => (x"87",x"c6",x"02",x"66"),
  1908 => (x"4a",x"d5",x"d5",x"c5"),
  1909 => (x"ff",x"cf",x"87",x"c4"),
  1910 => (x"e8",x"c2",x"4a",x"ff"),
  1911 => (x"e8",x"c2",x"5a",x"ce"),
  1912 => (x"78",x"c1",x"48",x"ce"),
  1913 => (x"26",x"87",x"c4",x"26"),
  1914 => (x"26",x"4c",x"26",x"4d"),
  1915 => (x"0e",x"4f",x"26",x"4b"),
  1916 => (x"5d",x"5c",x"5b",x"5e"),
  1917 => (x"c2",x"4a",x"71",x"0e"),
  1918 => (x"4c",x"bf",x"ca",x"e8"),
  1919 => (x"cb",x"02",x"9a",x"72"),
  1920 => (x"91",x"c8",x"49",x"87"),
  1921 => (x"4b",x"f0",x"f6",x"c1"),
  1922 => (x"87",x"c4",x"83",x"71"),
  1923 => (x"4b",x"f0",x"fa",x"c1"),
  1924 => (x"49",x"13",x"4d",x"c0"),
  1925 => (x"e8",x"c2",x"99",x"74"),
  1926 => (x"71",x"48",x"bf",x"c6"),
  1927 => (x"08",x"d4",x"ff",x"b8"),
  1928 => (x"2c",x"b7",x"c1",x"78"),
  1929 => (x"ad",x"b7",x"c8",x"85"),
  1930 => (x"c2",x"87",x"e7",x"04"),
  1931 => (x"48",x"bf",x"c2",x"e8"),
  1932 => (x"e8",x"c2",x"80",x"c8"),
  1933 => (x"ee",x"fe",x"58",x"c6"),
  1934 => (x"1e",x"73",x"1e",x"87"),
  1935 => (x"4a",x"13",x"4b",x"71"),
  1936 => (x"87",x"cb",x"02",x"9a"),
  1937 => (x"e6",x"fe",x"49",x"72"),
  1938 => (x"9a",x"4a",x"13",x"87"),
  1939 => (x"fe",x"87",x"f5",x"05"),
  1940 => (x"1e",x"1e",x"87",x"d9"),
  1941 => (x"bf",x"c2",x"e8",x"c2"),
  1942 => (x"c2",x"e8",x"c2",x"49"),
  1943 => (x"78",x"a1",x"c1",x"48"),
  1944 => (x"a9",x"b7",x"c0",x"c4"),
  1945 => (x"ff",x"87",x"db",x"03"),
  1946 => (x"e8",x"c2",x"48",x"d4"),
  1947 => (x"c2",x"78",x"bf",x"c6"),
  1948 => (x"49",x"bf",x"c2",x"e8"),
  1949 => (x"48",x"c2",x"e8",x"c2"),
  1950 => (x"c4",x"78",x"a1",x"c1"),
  1951 => (x"04",x"a9",x"b7",x"c0"),
  1952 => (x"d0",x"ff",x"87",x"e5"),
  1953 => (x"c0",x"c8",x"48",x"bf"),
  1954 => (x"a6",x"c4",x"98",x"c0"),
  1955 => (x"02",x"98",x"70",x"58"),
  1956 => (x"d0",x"ff",x"87",x"d0"),
  1957 => (x"c0",x"c8",x"48",x"bf"),
  1958 => (x"a6",x"c4",x"98",x"c0"),
  1959 => (x"05",x"98",x"70",x"58"),
  1960 => (x"d0",x"ff",x"87",x"f0"),
  1961 => (x"c2",x"78",x"c8",x"48"),
  1962 => (x"c0",x"48",x"ce",x"e8"),
  1963 => (x"4f",x"26",x"26",x"78"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"5f",x"00",x"00",x"00"),
  1967 => (x"00",x"00",x"00",x"5f"),
  1968 => (x"00",x"03",x"03",x"00"),
  1969 => (x"00",x"00",x"03",x"03"),
  1970 => (x"14",x"7f",x"7f",x"14"),
  1971 => (x"00",x"14",x"7f",x"7f"),
  1972 => (x"6b",x"2e",x"24",x"00"),
  1973 => (x"00",x"12",x"3a",x"6b"),
  1974 => (x"18",x"36",x"6a",x"4c"),
  1975 => (x"00",x"32",x"56",x"6c"),
  1976 => (x"59",x"4f",x"7e",x"30"),
  1977 => (x"40",x"68",x"3a",x"77"),
  1978 => (x"07",x"04",x"00",x"00"),
  1979 => (x"00",x"00",x"00",x"03"),
  1980 => (x"3e",x"1c",x"00",x"00"),
  1981 => (x"00",x"00",x"41",x"63"),
  1982 => (x"63",x"41",x"00",x"00"),
  1983 => (x"00",x"00",x"1c",x"3e"),
  1984 => (x"1c",x"3e",x"2a",x"08"),
  1985 => (x"08",x"2a",x"3e",x"1c"),
  1986 => (x"3e",x"08",x"08",x"00"),
  1987 => (x"00",x"08",x"08",x"3e"),
  1988 => (x"e0",x"80",x"00",x"00"),
  1989 => (x"00",x"00",x"00",x"60"),
  1990 => (x"08",x"08",x"08",x"00"),
  1991 => (x"00",x"08",x"08",x"08"),
  1992 => (x"60",x"00",x"00",x"00"),
  1993 => (x"00",x"00",x"00",x"60"),
  1994 => (x"18",x"30",x"60",x"40"),
  1995 => (x"01",x"03",x"06",x"0c"),
  1996 => (x"59",x"7f",x"3e",x"00"),
  1997 => (x"00",x"3e",x"7f",x"4d"),
  1998 => (x"7f",x"06",x"04",x"00"),
  1999 => (x"00",x"00",x"00",x"7f"),
  2000 => (x"71",x"63",x"42",x"00"),
  2001 => (x"00",x"46",x"4f",x"59"),
  2002 => (x"49",x"63",x"22",x"00"),
  2003 => (x"00",x"36",x"7f",x"49"),
  2004 => (x"13",x"16",x"1c",x"18"),
  2005 => (x"00",x"10",x"7f",x"7f"),
  2006 => (x"45",x"67",x"27",x"00"),
  2007 => (x"00",x"39",x"7d",x"45"),
  2008 => (x"4b",x"7e",x"3c",x"00"),
  2009 => (x"00",x"30",x"79",x"49"),
  2010 => (x"71",x"01",x"01",x"00"),
  2011 => (x"00",x"07",x"0f",x"79"),
  2012 => (x"49",x"7f",x"36",x"00"),
  2013 => (x"00",x"36",x"7f",x"49"),
  2014 => (x"49",x"4f",x"06",x"00"),
  2015 => (x"00",x"1e",x"3f",x"69"),
  2016 => (x"66",x"00",x"00",x"00"),
  2017 => (x"00",x"00",x"00",x"66"),
  2018 => (x"e6",x"80",x"00",x"00"),
  2019 => (x"00",x"00",x"00",x"66"),
  2020 => (x"14",x"08",x"08",x"00"),
  2021 => (x"00",x"22",x"22",x"14"),
  2022 => (x"14",x"14",x"14",x"00"),
  2023 => (x"00",x"14",x"14",x"14"),
  2024 => (x"14",x"22",x"22",x"00"),
  2025 => (x"00",x"08",x"08",x"14"),
  2026 => (x"51",x"03",x"02",x"00"),
  2027 => (x"00",x"06",x"0f",x"59"),
  2028 => (x"5d",x"41",x"7f",x"3e"),
  2029 => (x"00",x"1e",x"1f",x"55"),
  2030 => (x"09",x"7f",x"7e",x"00"),
  2031 => (x"00",x"7e",x"7f",x"09"),
  2032 => (x"49",x"7f",x"7f",x"00"),
  2033 => (x"00",x"36",x"7f",x"49"),
  2034 => (x"63",x"3e",x"1c",x"00"),
  2035 => (x"00",x"41",x"41",x"41"),
  2036 => (x"41",x"7f",x"7f",x"00"),
  2037 => (x"00",x"1c",x"3e",x"63"),
  2038 => (x"49",x"7f",x"7f",x"00"),
  2039 => (x"00",x"41",x"41",x"49"),
  2040 => (x"09",x"7f",x"7f",x"00"),
  2041 => (x"00",x"01",x"01",x"09"),
  2042 => (x"41",x"7f",x"3e",x"00"),
  2043 => (x"00",x"7a",x"7b",x"49"),
  2044 => (x"08",x"7f",x"7f",x"00"),
  2045 => (x"00",x"7f",x"7f",x"08"),
  2046 => (x"7f",x"41",x"00",x"00"),
  2047 => (x"00",x"00",x"41",x"7f"),
  2048 => (x"40",x"60",x"20",x"00"),
  2049 => (x"00",x"3f",x"7f",x"40"),
  2050 => (x"1c",x"08",x"7f",x"7f"),
  2051 => (x"00",x"41",x"63",x"36"),
  2052 => (x"40",x"7f",x"7f",x"00"),
  2053 => (x"00",x"40",x"40",x"40"),
  2054 => (x"0c",x"06",x"7f",x"7f"),
  2055 => (x"00",x"7f",x"7f",x"06"),
  2056 => (x"0c",x"06",x"7f",x"7f"),
  2057 => (x"00",x"7f",x"7f",x"18"),
  2058 => (x"41",x"7f",x"3e",x"00"),
  2059 => (x"00",x"3e",x"7f",x"41"),
  2060 => (x"09",x"7f",x"7f",x"00"),
  2061 => (x"00",x"06",x"0f",x"09"),
  2062 => (x"61",x"41",x"7f",x"3e"),
  2063 => (x"00",x"40",x"7e",x"7f"),
  2064 => (x"09",x"7f",x"7f",x"00"),
  2065 => (x"00",x"66",x"7f",x"19"),
  2066 => (x"4d",x"6f",x"26",x"00"),
  2067 => (x"00",x"32",x"7b",x"59"),
  2068 => (x"7f",x"01",x"01",x"00"),
  2069 => (x"00",x"01",x"01",x"7f"),
  2070 => (x"40",x"7f",x"3f",x"00"),
  2071 => (x"00",x"3f",x"7f",x"40"),
  2072 => (x"70",x"3f",x"0f",x"00"),
  2073 => (x"00",x"0f",x"3f",x"70"),
  2074 => (x"18",x"30",x"7f",x"7f"),
  2075 => (x"00",x"7f",x"7f",x"30"),
  2076 => (x"1c",x"36",x"63",x"41"),
  2077 => (x"41",x"63",x"36",x"1c"),
  2078 => (x"7c",x"06",x"03",x"01"),
  2079 => (x"01",x"03",x"06",x"7c"),
  2080 => (x"4d",x"59",x"71",x"61"),
  2081 => (x"00",x"41",x"43",x"47"),
  2082 => (x"7f",x"7f",x"00",x"00"),
  2083 => (x"00",x"00",x"41",x"41"),
  2084 => (x"0c",x"06",x"03",x"01"),
  2085 => (x"40",x"60",x"30",x"18"),
  2086 => (x"41",x"41",x"00",x"00"),
  2087 => (x"00",x"00",x"7f",x"7f"),
  2088 => (x"03",x"06",x"0c",x"08"),
  2089 => (x"00",x"08",x"0c",x"06"),
  2090 => (x"80",x"80",x"80",x"80"),
  2091 => (x"00",x"80",x"80",x"80"),
  2092 => (x"03",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"04",x"07"),
  2094 => (x"54",x"74",x"20",x"00"),
  2095 => (x"00",x"78",x"7c",x"54"),
  2096 => (x"44",x"7f",x"7f",x"00"),
  2097 => (x"00",x"38",x"7c",x"44"),
  2098 => (x"44",x"7c",x"38",x"00"),
  2099 => (x"00",x"00",x"44",x"44"),
  2100 => (x"44",x"7c",x"38",x"00"),
  2101 => (x"00",x"7f",x"7f",x"44"),
  2102 => (x"54",x"7c",x"38",x"00"),
  2103 => (x"00",x"18",x"5c",x"54"),
  2104 => (x"7f",x"7e",x"04",x"00"),
  2105 => (x"00",x"00",x"05",x"05"),
  2106 => (x"a4",x"bc",x"18",x"00"),
  2107 => (x"00",x"7c",x"fc",x"a4"),
  2108 => (x"04",x"7f",x"7f",x"00"),
  2109 => (x"00",x"78",x"7c",x"04"),
  2110 => (x"3d",x"00",x"00",x"00"),
  2111 => (x"00",x"00",x"40",x"7d"),
  2112 => (x"80",x"80",x"80",x"00"),
  2113 => (x"00",x"00",x"7d",x"fd"),
  2114 => (x"10",x"7f",x"7f",x"00"),
  2115 => (x"00",x"44",x"6c",x"38"),
  2116 => (x"3f",x"00",x"00",x"00"),
  2117 => (x"00",x"00",x"40",x"7f"),
  2118 => (x"18",x"0c",x"7c",x"7c"),
  2119 => (x"00",x"78",x"7c",x"0c"),
  2120 => (x"04",x"7c",x"7c",x"00"),
  2121 => (x"00",x"78",x"7c",x"04"),
  2122 => (x"44",x"7c",x"38",x"00"),
  2123 => (x"00",x"38",x"7c",x"44"),
  2124 => (x"24",x"fc",x"fc",x"00"),
  2125 => (x"00",x"18",x"3c",x"24"),
  2126 => (x"24",x"3c",x"18",x"00"),
  2127 => (x"00",x"fc",x"fc",x"24"),
  2128 => (x"04",x"7c",x"7c",x"00"),
  2129 => (x"00",x"08",x"0c",x"04"),
  2130 => (x"54",x"5c",x"48",x"00"),
  2131 => (x"00",x"20",x"74",x"54"),
  2132 => (x"7f",x"3f",x"04",x"00"),
  2133 => (x"00",x"00",x"44",x"44"),
  2134 => (x"40",x"7c",x"3c",x"00"),
  2135 => (x"00",x"7c",x"7c",x"40"),
  2136 => (x"60",x"3c",x"1c",x"00"),
  2137 => (x"00",x"1c",x"3c",x"60"),
  2138 => (x"30",x"60",x"7c",x"3c"),
  2139 => (x"00",x"3c",x"7c",x"60"),
  2140 => (x"10",x"38",x"6c",x"44"),
  2141 => (x"00",x"44",x"6c",x"38"),
  2142 => (x"e0",x"bc",x"1c",x"00"),
  2143 => (x"00",x"1c",x"3c",x"60"),
  2144 => (x"74",x"64",x"44",x"00"),
  2145 => (x"00",x"44",x"4c",x"5c"),
  2146 => (x"3e",x"08",x"08",x"00"),
  2147 => (x"00",x"41",x"41",x"77"),
  2148 => (x"7f",x"00",x"00",x"00"),
  2149 => (x"00",x"00",x"00",x"7f"),
  2150 => (x"77",x"41",x"41",x"00"),
  2151 => (x"00",x"08",x"08",x"3e"),
  2152 => (x"03",x"01",x"01",x"02"),
  2153 => (x"00",x"01",x"02",x"02"),
  2154 => (x"7f",x"7f",x"7f",x"7f"),
  2155 => (x"00",x"7f",x"7f",x"7f"),
  2156 => (x"1c",x"1c",x"08",x"08"),
  2157 => (x"7f",x"7f",x"3e",x"3e"),
  2158 => (x"3e",x"3e",x"7f",x"7f"),
  2159 => (x"08",x"08",x"1c",x"1c"),
  2160 => (x"7c",x"18",x"10",x"00"),
  2161 => (x"00",x"10",x"18",x"7c"),
  2162 => (x"7c",x"30",x"10",x"00"),
  2163 => (x"00",x"10",x"30",x"7c"),
  2164 => (x"60",x"60",x"30",x"10"),
  2165 => (x"00",x"06",x"1e",x"78"),
  2166 => (x"18",x"3c",x"66",x"42"),
  2167 => (x"00",x"42",x"66",x"3c"),
  2168 => (x"c2",x"6a",x"38",x"78"),
  2169 => (x"00",x"38",x"6c",x"c6"),
  2170 => (x"60",x"00",x"00",x"60"),
  2171 => (x"00",x"60",x"00",x"00"),
  2172 => (x"5c",x"5b",x"5e",x"0e"),
  2173 => (x"71",x"1e",x"0e",x"5d"),
  2174 => (x"d6",x"e8",x"c2",x"4c"),
  2175 => (x"4b",x"c0",x"4d",x"bf"),
  2176 => (x"ab",x"74",x"1e",x"c0"),
  2177 => (x"c4",x"87",x"c7",x"02"),
  2178 => (x"78",x"c0",x"48",x"a6"),
  2179 => (x"a6",x"c4",x"87",x"c5"),
  2180 => (x"c4",x"78",x"c1",x"48"),
  2181 => (x"49",x"73",x"1e",x"66"),
  2182 => (x"c8",x"87",x"db",x"ed"),
  2183 => (x"49",x"e0",x"c0",x"86"),
  2184 => (x"c4",x"87",x"cc",x"ef"),
  2185 => (x"49",x"6a",x"4a",x"a5"),
  2186 => (x"f0",x"87",x"ce",x"f0"),
  2187 => (x"85",x"cb",x"87",x"e4"),
  2188 => (x"b7",x"c8",x"83",x"c1"),
  2189 => (x"c7",x"ff",x"04",x"ab"),
  2190 => (x"4d",x"26",x"26",x"87"),
  2191 => (x"4b",x"26",x"4c",x"26"),
  2192 => (x"71",x"1e",x"4f",x"26"),
  2193 => (x"da",x"e8",x"c2",x"4a"),
  2194 => (x"da",x"e8",x"c2",x"5a"),
  2195 => (x"49",x"78",x"c7",x"48"),
  2196 => (x"26",x"87",x"dd",x"fe"),
  2197 => (x"c0",x"c1",x"1e",x"4f"),
  2198 => (x"87",x"ea",x"eb",x"49"),
  2199 => (x"48",x"c5",x"d3",x"c2"),
  2200 => (x"4f",x"26",x"78",x"c0"),
  2201 => (x"5c",x"5b",x"5e",x"0e"),
  2202 => (x"86",x"f4",x"0e",x"5d"),
  2203 => (x"a6",x"c8",x"7e",x"c0"),
  2204 => (x"78",x"bf",x"ec",x"48"),
  2205 => (x"e8",x"c2",x"80",x"fc"),
  2206 => (x"c2",x"78",x"bf",x"d6"),
  2207 => (x"4d",x"bf",x"de",x"e8"),
  2208 => (x"c7",x"4c",x"bf",x"e8"),
  2209 => (x"87",x"c9",x"e7",x"49"),
  2210 => (x"99",x"c2",x"49",x"70"),
  2211 => (x"c2",x"87",x"d0",x"05"),
  2212 => (x"49",x"bf",x"fd",x"d2"),
  2213 => (x"66",x"c8",x"b9",x"ff"),
  2214 => (x"02",x"99",x"c1",x"99"),
  2215 => (x"c7",x"87",x"eb",x"c0"),
  2216 => (x"87",x"ed",x"e6",x"49"),
  2217 => (x"cd",x"02",x"98",x"70"),
  2218 => (x"87",x"db",x"e2",x"87"),
  2219 => (x"e0",x"e6",x"49",x"c7"),
  2220 => (x"05",x"98",x"70",x"87"),
  2221 => (x"d3",x"c2",x"87",x"f3"),
  2222 => (x"c1",x"4a",x"bf",x"c5"),
  2223 => (x"c9",x"d3",x"c2",x"ba"),
  2224 => (x"a2",x"c0",x"c1",x"5a"),
  2225 => (x"87",x"fe",x"e9",x"49"),
  2226 => (x"d2",x"c2",x"7e",x"c1"),
  2227 => (x"66",x"c8",x"48",x"fd"),
  2228 => (x"c5",x"d3",x"c2",x"78"),
  2229 => (x"cb",x"c1",x"05",x"bf"),
  2230 => (x"c0",x"c0",x"c8",x"87"),
  2231 => (x"c9",x"d3",x"c2",x"7e"),
  2232 => (x"e5",x"49",x"13",x"4b"),
  2233 => (x"98",x"70",x"87",x"eb"),
  2234 => (x"6e",x"87",x"c2",x"02"),
  2235 => (x"c1",x"48",x"6e",x"b4"),
  2236 => (x"a6",x"c4",x"28",x"b7"),
  2237 => (x"05",x"98",x"70",x"58"),
  2238 => (x"74",x"87",x"e6",x"ff"),
  2239 => (x"99",x"ff",x"c3",x"49"),
  2240 => (x"49",x"c0",x"1e",x"71"),
  2241 => (x"74",x"87",x"f2",x"e7"),
  2242 => (x"29",x"b7",x"c8",x"49"),
  2243 => (x"49",x"c1",x"1e",x"71"),
  2244 => (x"c8",x"87",x"e6",x"e7"),
  2245 => (x"49",x"fd",x"c3",x"86"),
  2246 => (x"c3",x"87",x"f6",x"e4"),
  2247 => (x"f0",x"e4",x"49",x"fa"),
  2248 => (x"87",x"c4",x"c6",x"87"),
  2249 => (x"ff",x"c3",x"49",x"74"),
  2250 => (x"2c",x"b7",x"c8",x"99"),
  2251 => (x"9c",x"74",x"b4",x"71"),
  2252 => (x"87",x"e2",x"c0",x"02"),
  2253 => (x"ff",x"48",x"a6",x"c8"),
  2254 => (x"c8",x"78",x"bf",x"c8"),
  2255 => (x"d3",x"c2",x"49",x"66"),
  2256 => (x"c2",x"89",x"bf",x"c1"),
  2257 => (x"c4",x"03",x"a9",x"e0"),
  2258 => (x"cf",x"4c",x"c0",x"87"),
  2259 => (x"c1",x"d3",x"c2",x"87"),
  2260 => (x"78",x"66",x"c8",x"48"),
  2261 => (x"d3",x"c2",x"87",x"c6"),
  2262 => (x"78",x"c0",x"48",x"c1"),
  2263 => (x"99",x"c8",x"49",x"74"),
  2264 => (x"c3",x"87",x"ce",x"05"),
  2265 => (x"e8",x"e3",x"49",x"f5"),
  2266 => (x"c2",x"49",x"70",x"87"),
  2267 => (x"e6",x"c0",x"02",x"99"),
  2268 => (x"da",x"e8",x"c2",x"87"),
  2269 => (x"87",x"c9",x"02",x"bf"),
  2270 => (x"c2",x"88",x"c1",x"48"),
  2271 => (x"d4",x"58",x"de",x"e8"),
  2272 => (x"48",x"66",x"c4",x"87"),
  2273 => (x"c4",x"80",x"d8",x"c1"),
  2274 => (x"bf",x"6e",x"58",x"a6"),
  2275 => (x"87",x"c5",x"c0",x"02"),
  2276 => (x"73",x"49",x"ff",x"4b"),
  2277 => (x"74",x"7e",x"c1",x"0f"),
  2278 => (x"05",x"99",x"c4",x"49"),
  2279 => (x"f2",x"c3",x"87",x"ce"),
  2280 => (x"87",x"ed",x"e2",x"49"),
  2281 => (x"99",x"c2",x"49",x"70"),
  2282 => (x"87",x"ee",x"c0",x"02"),
  2283 => (x"bf",x"da",x"e8",x"c2"),
  2284 => (x"c7",x"48",x"6e",x"7e"),
  2285 => (x"c0",x"03",x"a8",x"b7"),
  2286 => (x"48",x"6e",x"87",x"ca"),
  2287 => (x"e8",x"c2",x"80",x"c1"),
  2288 => (x"87",x"d4",x"58",x"de"),
  2289 => (x"c1",x"48",x"66",x"c4"),
  2290 => (x"a6",x"c4",x"80",x"d8"),
  2291 => (x"02",x"bf",x"6e",x"58"),
  2292 => (x"4b",x"87",x"c5",x"c0"),
  2293 => (x"0f",x"73",x"49",x"fe"),
  2294 => (x"fd",x"c3",x"7e",x"c1"),
  2295 => (x"87",x"f1",x"e1",x"49"),
  2296 => (x"99",x"c2",x"49",x"70"),
  2297 => (x"87",x"e3",x"c0",x"02"),
  2298 => (x"bf",x"da",x"e8",x"c2"),
  2299 => (x"87",x"c9",x"c0",x"02"),
  2300 => (x"48",x"da",x"e8",x"c2"),
  2301 => (x"d0",x"c0",x"78",x"c0"),
  2302 => (x"4a",x"66",x"c4",x"87"),
  2303 => (x"6a",x"82",x"d8",x"c1"),
  2304 => (x"87",x"c5",x"c0",x"02"),
  2305 => (x"73",x"49",x"fd",x"4b"),
  2306 => (x"c3",x"7e",x"c1",x"0f"),
  2307 => (x"c0",x"e1",x"49",x"fa"),
  2308 => (x"c2",x"49",x"70",x"87"),
  2309 => (x"eb",x"c0",x"02",x"99"),
  2310 => (x"da",x"e8",x"c2",x"87"),
  2311 => (x"b7",x"c7",x"48",x"bf"),
  2312 => (x"c9",x"c0",x"03",x"a8"),
  2313 => (x"da",x"e8",x"c2",x"87"),
  2314 => (x"c0",x"78",x"c7",x"48"),
  2315 => (x"66",x"c4",x"87",x"d4"),
  2316 => (x"80",x"d8",x"c1",x"48"),
  2317 => (x"6e",x"58",x"a6",x"c4"),
  2318 => (x"c5",x"c0",x"02",x"bf"),
  2319 => (x"49",x"fc",x"4b",x"87"),
  2320 => (x"7e",x"c1",x"0f",x"73"),
  2321 => (x"f0",x"c3",x"49",x"74"),
  2322 => (x"cf",x"c0",x"05",x"99"),
  2323 => (x"49",x"da",x"c1",x"87"),
  2324 => (x"87",x"fd",x"df",x"ff"),
  2325 => (x"99",x"c2",x"49",x"70"),
  2326 => (x"87",x"d0",x"c0",x"02"),
  2327 => (x"bf",x"da",x"e8",x"c2"),
  2328 => (x"93",x"cb",x"4b",x"49"),
  2329 => (x"6b",x"83",x"66",x"c4"),
  2330 => (x"0f",x"73",x"71",x"4b"),
  2331 => (x"c0",x"02",x"9d",x"75"),
  2332 => (x"02",x"6d",x"87",x"e9"),
  2333 => (x"6d",x"87",x"e4",x"c0"),
  2334 => (x"d4",x"df",x"ff",x"49"),
  2335 => (x"c1",x"49",x"70",x"87"),
  2336 => (x"cb",x"c0",x"02",x"99"),
  2337 => (x"4b",x"a5",x"c4",x"87"),
  2338 => (x"bf",x"da",x"e8",x"c2"),
  2339 => (x"0f",x"4b",x"6b",x"49"),
  2340 => (x"c0",x"02",x"85",x"c8"),
  2341 => (x"05",x"6d",x"87",x"c5"),
  2342 => (x"6e",x"87",x"dc",x"ff"),
  2343 => (x"87",x"c8",x"c0",x"02"),
  2344 => (x"bf",x"da",x"e8",x"c2"),
  2345 => (x"87",x"c8",x"f5",x"49"),
  2346 => (x"cd",x"f6",x"8e",x"f4"),
  2347 => (x"11",x"12",x"58",x"87"),
  2348 => (x"1c",x"1b",x"1d",x"14"),
  2349 => (x"91",x"59",x"5a",x"23"),
  2350 => (x"eb",x"f2",x"f5",x"94"),
  2351 => (x"00",x"00",x"00",x"f4"),
  2352 => (x"00",x"00",x"00",x"00"),
  2353 => (x"00",x"00",x"00",x"00"),
  2354 => (x"14",x"12",x"58",x"00"),
  2355 => (x"1c",x"1b",x"1d",x"11"),
  2356 => (x"94",x"59",x"5a",x"23"),
  2357 => (x"eb",x"f2",x"f5",x"91"),
  2358 => (x"00",x"00",x"00",x"f4"),
  2359 => (x"00",x"00",x"24",x"e0"),
  2360 => (x"4f",x"54",x"55",x"41"),
  2361 => (x"54",x"4f",x"4f",x"42"),
  2362 => (x"00",x"53",x"45",x"4e"),
  2363 => (x"00",x"00",x"19",x"c6"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

