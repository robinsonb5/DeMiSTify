
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"ec",x"c2",x"87"),
    12 => (x"48",x"c0",x"c4",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"05",x"88"),
    17 => (x"49",x"d8",x"ec",x"c2"),
    18 => (x"48",x"e4",x"d7",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"e4",x"d7",x"c2",x"87"),
    25 => (x"e0",x"d7",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e1",x"c1",x"87",x"f7"),
    29 => (x"d7",x"c2",x"87",x"c1"),
    30 => (x"d7",x"c2",x"4d",x"e4"),
    31 => (x"ad",x"74",x"4c",x"e4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"c0",x"4b",x"71",x"0e"),
    37 => (x"9a",x"4a",x"13",x"4c"),
    38 => (x"72",x"87",x"cd",x"02"),
    39 => (x"87",x"e0",x"c0",x"49"),
    40 => (x"4a",x"13",x"84",x"c1"),
    41 => (x"87",x"f3",x"05",x"9a"),
    42 => (x"4c",x"26",x"48",x"74"),
    43 => (x"4f",x"26",x"4b",x"26"),
    44 => (x"81",x"48",x"73",x"1e"),
    45 => (x"c5",x"02",x"a9",x"73"),
    46 => (x"05",x"53",x"12",x"87"),
    47 => (x"4f",x"26",x"87",x"f6"),
    48 => (x"c0",x"ff",x"1e",x"1e"),
    49 => (x"c4",x"48",x"6a",x"4a"),
    50 => (x"a6",x"c4",x"98",x"c0"),
    51 => (x"02",x"98",x"70",x"58"),
    52 => (x"7a",x"71",x"87",x"f3"),
    53 => (x"4f",x"26",x"26",x"48"),
    54 => (x"ff",x"1e",x"73",x"1e"),
    55 => (x"ff",x"c3",x"4b",x"d4"),
    56 => (x"c3",x"4a",x"6b",x"7b"),
    57 => (x"49",x"6b",x"7b",x"ff"),
    58 => (x"b1",x"72",x"32",x"c8"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"71",x"31",x"c8",x"4a"),
    61 => (x"7b",x"ff",x"c3",x"b2"),
    62 => (x"32",x"c8",x"49",x"6b"),
    63 => (x"48",x"71",x"b1",x"72"),
    64 => (x"4d",x"26",x"87",x"c4"),
    65 => (x"4b",x"26",x"4c",x"26"),
    66 => (x"5e",x"0e",x"4f",x"26"),
    67 => (x"0e",x"5d",x"5c",x"5b"),
    68 => (x"d4",x"ff",x"4a",x"71"),
    69 => (x"c3",x"48",x"72",x"4c"),
    70 => (x"7c",x"70",x"98",x"ff"),
    71 => (x"bf",x"e4",x"d7",x"c2"),
    72 => (x"d0",x"87",x"c8",x"05"),
    73 => (x"30",x"c9",x"48",x"66"),
    74 => (x"d0",x"58",x"a6",x"d4"),
    75 => (x"29",x"d8",x"49",x"66"),
    76 => (x"ff",x"c3",x"48",x"71"),
    77 => (x"d0",x"7c",x"70",x"98"),
    78 => (x"29",x"d0",x"49",x"66"),
    79 => (x"ff",x"c3",x"48",x"71"),
    80 => (x"d0",x"7c",x"70",x"98"),
    81 => (x"29",x"c8",x"49",x"66"),
    82 => (x"ff",x"c3",x"48",x"71"),
    83 => (x"d0",x"7c",x"70",x"98"),
    84 => (x"ff",x"c3",x"48",x"66"),
    85 => (x"72",x"7c",x"70",x"98"),
    86 => (x"71",x"29",x"d0",x"49"),
    87 => (x"98",x"ff",x"c3",x"48"),
    88 => (x"4b",x"6c",x"7c",x"70"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"ff",x"fd"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"df",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c1",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"de",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"49",x"e3",x"c8",x"78"),
   125 => (x"d3",x"87",x"d5",x"fa"),
   126 => (x"c0",x"1e",x"c0",x"4b"),
   127 => (x"c1",x"c1",x"f0",x"ff"),
   128 => (x"87",x"c6",x"fc",x"49"),
   129 => (x"98",x"70",x"86",x"c4"),
   130 => (x"ff",x"87",x"ca",x"05"),
   131 => (x"ff",x"c3",x"48",x"d4"),
   132 => (x"cb",x"48",x"c1",x"78"),
   133 => (x"87",x"eb",x"fd",x"87"),
   134 => (x"ff",x"05",x"8b",x"c1"),
   135 => (x"48",x"c0",x"87",x"db"),
   136 => (x"43",x"87",x"e3",x"fb"),
   137 => (x"53",x"00",x"44",x"4d"),
   138 => (x"20",x"43",x"48",x"44"),
   139 => (x"6c",x"69",x"61",x"66"),
   140 => (x"49",x"00",x"0a",x"21"),
   141 => (x"00",x"52",x"52",x"45"),
   142 => (x"00",x"49",x"50",x"53"),
   143 => (x"74",x"69",x"72",x"57"),
   144 => (x"61",x"66",x"20",x"65"),
   145 => (x"64",x"65",x"6c",x"69"),
   146 => (x"5e",x"0e",x"00",x"0a"),
   147 => (x"ff",x"0e",x"5c",x"5b"),
   148 => (x"ee",x"fc",x"4c",x"d4"),
   149 => (x"1e",x"ea",x"c6",x"87"),
   150 => (x"c1",x"f0",x"e1",x"c0"),
   151 => (x"e9",x"fa",x"49",x"c8"),
   152 => (x"c1",x"86",x"c4",x"87"),
   153 => (x"87",x"c8",x"02",x"a8"),
   154 => (x"c0",x"87",x"fd",x"fd"),
   155 => (x"87",x"e8",x"c1",x"48"),
   156 => (x"70",x"87",x"e5",x"f9"),
   157 => (x"ff",x"ff",x"cf",x"49"),
   158 => (x"a9",x"ea",x"c6",x"99"),
   159 => (x"fd",x"87",x"c8",x"02"),
   160 => (x"48",x"c0",x"87",x"e6"),
   161 => (x"c3",x"87",x"d1",x"c1"),
   162 => (x"f1",x"c0",x"7c",x"ff"),
   163 => (x"87",x"c7",x"fc",x"4b"),
   164 => (x"c0",x"02",x"98",x"70"),
   165 => (x"1e",x"c0",x"87",x"eb"),
   166 => (x"c1",x"f0",x"ff",x"c0"),
   167 => (x"e9",x"f9",x"49",x"fa"),
   168 => (x"70",x"86",x"c4",x"87"),
   169 => (x"87",x"d9",x"05",x"98"),
   170 => (x"6c",x"7c",x"ff",x"c3"),
   171 => (x"7c",x"ff",x"c3",x"49"),
   172 => (x"c1",x"7c",x"7c",x"7c"),
   173 => (x"c4",x"02",x"99",x"c0"),
   174 => (x"db",x"48",x"c1",x"87"),
   175 => (x"d7",x"48",x"c0",x"87"),
   176 => (x"05",x"ab",x"c2",x"87"),
   177 => (x"e7",x"c8",x"87",x"ca"),
   178 => (x"87",x"c0",x"f7",x"49"),
   179 => (x"87",x"c8",x"48",x"c0"),
   180 => (x"fe",x"05",x"8b",x"c1"),
   181 => (x"48",x"c0",x"87",x"f7"),
   182 => (x"0e",x"87",x"e9",x"f8"),
   183 => (x"5d",x"5c",x"5b",x"5e"),
   184 => (x"d0",x"ff",x"1e",x"0e"),
   185 => (x"c0",x"c0",x"c8",x"4d"),
   186 => (x"e4",x"d7",x"c2",x"4b"),
   187 => (x"c8",x"78",x"c1",x"48"),
   188 => (x"d7",x"f6",x"49",x"f8"),
   189 => (x"6d",x"4c",x"c7",x"87"),
   190 => (x"c4",x"98",x"73",x"48"),
   191 => (x"98",x"70",x"58",x"a6"),
   192 => (x"6d",x"87",x"cc",x"02"),
   193 => (x"c4",x"98",x"73",x"48"),
   194 => (x"98",x"70",x"58",x"a6"),
   195 => (x"c2",x"87",x"f4",x"05"),
   196 => (x"87",x"ef",x"f9",x"7d"),
   197 => (x"98",x"73",x"48",x"6d"),
   198 => (x"70",x"58",x"a6",x"c4"),
   199 => (x"87",x"cc",x"02",x"98"),
   200 => (x"98",x"73",x"48",x"6d"),
   201 => (x"70",x"58",x"a6",x"c4"),
   202 => (x"87",x"f4",x"05",x"98"),
   203 => (x"1e",x"c0",x"7d",x"c3"),
   204 => (x"c1",x"d0",x"e5",x"c0"),
   205 => (x"d1",x"f7",x"49",x"c0"),
   206 => (x"c1",x"86",x"c4",x"87"),
   207 => (x"87",x"c1",x"05",x"a8"),
   208 => (x"05",x"ac",x"c2",x"4c"),
   209 => (x"f3",x"c8",x"87",x"cb"),
   210 => (x"87",x"c0",x"f5",x"49"),
   211 => (x"ce",x"c1",x"48",x"c0"),
   212 => (x"05",x"8c",x"c1",x"87"),
   213 => (x"fb",x"87",x"e0",x"fe"),
   214 => (x"d7",x"c2",x"87",x"f0"),
   215 => (x"98",x"70",x"58",x"e8"),
   216 => (x"c1",x"87",x"cd",x"05"),
   217 => (x"f0",x"ff",x"c0",x"1e"),
   218 => (x"f6",x"49",x"d0",x"c1"),
   219 => (x"86",x"c4",x"87",x"dc"),
   220 => (x"c3",x"48",x"d4",x"ff"),
   221 => (x"dd",x"c5",x"78",x"ff"),
   222 => (x"ec",x"d7",x"c2",x"87"),
   223 => (x"73",x"48",x"6d",x"58"),
   224 => (x"58",x"a6",x"c4",x"98"),
   225 => (x"cc",x"02",x"98",x"70"),
   226 => (x"73",x"48",x"6d",x"87"),
   227 => (x"58",x"a6",x"c4",x"98"),
   228 => (x"f4",x"05",x"98",x"70"),
   229 => (x"ff",x"7d",x"c2",x"87"),
   230 => (x"ff",x"c3",x"48",x"d4"),
   231 => (x"26",x"48",x"c1",x"78"),
   232 => (x"0e",x"87",x"df",x"f5"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"c8",x"1e",x"0e"),
   235 => (x"4c",x"c0",x"4b",x"c0"),
   236 => (x"df",x"cd",x"ee",x"c5"),
   237 => (x"5c",x"a6",x"c4",x"4a"),
   238 => (x"c3",x"4c",x"d4",x"ff"),
   239 => (x"48",x"6c",x"7c",x"ff"),
   240 => (x"05",x"a8",x"fe",x"c3"),
   241 => (x"71",x"87",x"c0",x"c2"),
   242 => (x"e2",x"c0",x"05",x"99"),
   243 => (x"bf",x"d0",x"ff",x"87"),
   244 => (x"c4",x"98",x"73",x"48"),
   245 => (x"98",x"70",x"58",x"a6"),
   246 => (x"ff",x"87",x"ce",x"02"),
   247 => (x"73",x"48",x"bf",x"d0"),
   248 => (x"58",x"a6",x"c4",x"98"),
   249 => (x"f2",x"05",x"98",x"70"),
   250 => (x"48",x"d0",x"ff",x"87"),
   251 => (x"d4",x"78",x"d1",x"c4"),
   252 => (x"b7",x"c0",x"48",x"66"),
   253 => (x"e0",x"c0",x"06",x"a8"),
   254 => (x"7c",x"ff",x"c3",x"87"),
   255 => (x"99",x"71",x"4a",x"6c"),
   256 => (x"71",x"87",x"c7",x"02"),
   257 => (x"0a",x"7a",x"97",x"0a"),
   258 => (x"66",x"d4",x"81",x"c1"),
   259 => (x"d8",x"88",x"c1",x"48"),
   260 => (x"b7",x"c0",x"58",x"a6"),
   261 => (x"e0",x"ff",x"01",x"a8"),
   262 => (x"7c",x"ff",x"c3",x"87"),
   263 => (x"05",x"99",x"71",x"7c"),
   264 => (x"ff",x"87",x"e1",x"c0"),
   265 => (x"73",x"48",x"bf",x"d0"),
   266 => (x"58",x"a6",x"c4",x"98"),
   267 => (x"ce",x"02",x"98",x"70"),
   268 => (x"bf",x"d0",x"ff",x"87"),
   269 => (x"c4",x"98",x"73",x"48"),
   270 => (x"98",x"70",x"58",x"a6"),
   271 => (x"ff",x"87",x"f2",x"05"),
   272 => (x"78",x"d0",x"48",x"d0"),
   273 => (x"c1",x"7e",x"4a",x"c1"),
   274 => (x"ee",x"fd",x"05",x"8a"),
   275 => (x"26",x"48",x"6e",x"87"),
   276 => (x"0e",x"87",x"ef",x"f2"),
   277 => (x"0e",x"5c",x"5b",x"5e"),
   278 => (x"c8",x"4a",x"71",x"1e"),
   279 => (x"c0",x"4b",x"c0",x"c0"),
   280 => (x"48",x"d4",x"ff",x"4c"),
   281 => (x"ff",x"78",x"ff",x"c3"),
   282 => (x"73",x"48",x"bf",x"d0"),
   283 => (x"58",x"a6",x"c4",x"98"),
   284 => (x"ce",x"02",x"98",x"70"),
   285 => (x"bf",x"d0",x"ff",x"87"),
   286 => (x"c4",x"98",x"73",x"48"),
   287 => (x"98",x"70",x"58",x"a6"),
   288 => (x"ff",x"87",x"f2",x"05"),
   289 => (x"c3",x"c4",x"48",x"d0"),
   290 => (x"48",x"d4",x"ff",x"78"),
   291 => (x"72",x"78",x"ff",x"c3"),
   292 => (x"f0",x"ff",x"c0",x"1e"),
   293 => (x"f1",x"49",x"d1",x"c1"),
   294 => (x"86",x"c4",x"87",x"f0"),
   295 => (x"c0",x"05",x"98",x"70"),
   296 => (x"c0",x"c8",x"87",x"ee"),
   297 => (x"49",x"66",x"d4",x"1e"),
   298 => (x"c4",x"87",x"f8",x"fb"),
   299 => (x"ff",x"4c",x"70",x"86"),
   300 => (x"73",x"48",x"bf",x"d0"),
   301 => (x"58",x"a6",x"c4",x"98"),
   302 => (x"ce",x"02",x"98",x"70"),
   303 => (x"bf",x"d0",x"ff",x"87"),
   304 => (x"c4",x"98",x"73",x"48"),
   305 => (x"98",x"70",x"58",x"a6"),
   306 => (x"ff",x"87",x"f2",x"05"),
   307 => (x"78",x"c2",x"48",x"d0"),
   308 => (x"f0",x"26",x"48",x"74"),
   309 => (x"5e",x"0e",x"87",x"ee"),
   310 => (x"0e",x"5d",x"5c",x"5b"),
   311 => (x"ff",x"c0",x"1e",x"c0"),
   312 => (x"49",x"c9",x"c1",x"f0"),
   313 => (x"d2",x"87",x"e3",x"f0"),
   314 => (x"f2",x"d7",x"c2",x"1e"),
   315 => (x"87",x"f3",x"fa",x"49"),
   316 => (x"4c",x"c0",x"86",x"c8"),
   317 => (x"b7",x"d2",x"84",x"c1"),
   318 => (x"87",x"f8",x"04",x"ac"),
   319 => (x"97",x"f2",x"d7",x"c2"),
   320 => (x"c0",x"c3",x"49",x"bf"),
   321 => (x"a9",x"c0",x"c1",x"99"),
   322 => (x"87",x"e7",x"c0",x"05"),
   323 => (x"97",x"f9",x"d7",x"c2"),
   324 => (x"31",x"d0",x"49",x"bf"),
   325 => (x"97",x"fa",x"d7",x"c2"),
   326 => (x"32",x"c8",x"4a",x"bf"),
   327 => (x"d7",x"c2",x"b1",x"72"),
   328 => (x"4a",x"bf",x"97",x"fb"),
   329 => (x"cf",x"4c",x"71",x"b1"),
   330 => (x"9c",x"ff",x"ff",x"ff"),
   331 => (x"34",x"ca",x"84",x"c1"),
   332 => (x"c2",x"87",x"e7",x"c1"),
   333 => (x"bf",x"97",x"fb",x"d7"),
   334 => (x"c6",x"31",x"c1",x"49"),
   335 => (x"fc",x"d7",x"c2",x"99"),
   336 => (x"c7",x"4a",x"bf",x"97"),
   337 => (x"b1",x"72",x"2a",x"b7"),
   338 => (x"97",x"f7",x"d7",x"c2"),
   339 => (x"cf",x"4d",x"4a",x"bf"),
   340 => (x"f8",x"d7",x"c2",x"9d"),
   341 => (x"c3",x"4a",x"bf",x"97"),
   342 => (x"c2",x"32",x"ca",x"9a"),
   343 => (x"bf",x"97",x"f9",x"d7"),
   344 => (x"73",x"33",x"c2",x"4b"),
   345 => (x"fa",x"d7",x"c2",x"b2"),
   346 => (x"c3",x"4b",x"bf",x"97"),
   347 => (x"b7",x"c6",x"9b",x"c0"),
   348 => (x"c2",x"b2",x"73",x"2b"),
   349 => (x"71",x"48",x"c1",x"81"),
   350 => (x"c1",x"49",x"70",x"30"),
   351 => (x"70",x"30",x"75",x"48"),
   352 => (x"c1",x"4c",x"72",x"4d"),
   353 => (x"c8",x"94",x"71",x"84"),
   354 => (x"06",x"ad",x"b7",x"c0"),
   355 => (x"34",x"c1",x"87",x"cc"),
   356 => (x"c0",x"c8",x"2d",x"b7"),
   357 => (x"ff",x"01",x"ad",x"b7"),
   358 => (x"48",x"74",x"87",x"f4"),
   359 => (x"0e",x"87",x"e3",x"ed"),
   360 => (x"0e",x"5c",x"5b",x"5e"),
   361 => (x"4c",x"c0",x"4b",x"71"),
   362 => (x"c0",x"48",x"66",x"d0"),
   363 => (x"c0",x"06",x"a8",x"b7"),
   364 => (x"4a",x"13",x"87",x"e3"),
   365 => (x"bf",x"97",x"66",x"cc"),
   366 => (x"48",x"66",x"cc",x"49"),
   367 => (x"a6",x"d0",x"80",x"c1"),
   368 => (x"aa",x"b7",x"71",x"58"),
   369 => (x"c1",x"87",x"c4",x"02"),
   370 => (x"c1",x"87",x"cc",x"48"),
   371 => (x"b7",x"66",x"d0",x"84"),
   372 => (x"dd",x"ff",x"04",x"ac"),
   373 => (x"c2",x"48",x"c0",x"87"),
   374 => (x"26",x"4d",x"26",x"87"),
   375 => (x"26",x"4b",x"26",x"4c"),
   376 => (x"5b",x"5e",x"0e",x"4f"),
   377 => (x"c2",x"0e",x"5d",x"5c"),
   378 => (x"c0",x"48",x"d8",x"e0"),
   379 => (x"d0",x"d8",x"c2",x"78"),
   380 => (x"f9",x"49",x"c0",x"1e"),
   381 => (x"86",x"c4",x"87",x"dd"),
   382 => (x"c5",x"05",x"98",x"70"),
   383 => (x"c8",x"48",x"c0",x"87"),
   384 => (x"4b",x"c0",x"87",x"ef"),
   385 => (x"48",x"d0",x"e5",x"c2"),
   386 => (x"1e",x"c8",x"78",x"c1"),
   387 => (x"1e",x"fd",x"e0",x"c0"),
   388 => (x"49",x"c6",x"d9",x"c2"),
   389 => (x"c8",x"87",x"c8",x"fe"),
   390 => (x"05",x"98",x"70",x"86"),
   391 => (x"e5",x"c2",x"87",x"c6"),
   392 => (x"78",x"c0",x"48",x"d0"),
   393 => (x"e1",x"c0",x"1e",x"c8"),
   394 => (x"d9",x"c2",x"1e",x"c6"),
   395 => (x"ee",x"fd",x"49",x"e2"),
   396 => (x"70",x"86",x"c8",x"87"),
   397 => (x"87",x"c6",x"05",x"98"),
   398 => (x"48",x"d0",x"e5",x"c2"),
   399 => (x"e5",x"c2",x"78",x"c0"),
   400 => (x"c0",x"02",x"bf",x"d0"),
   401 => (x"df",x"c2",x"87",x"fa"),
   402 => (x"c2",x"4b",x"bf",x"d6"),
   403 => (x"bf",x"9f",x"ce",x"e0"),
   404 => (x"ea",x"d6",x"c5",x"4a"),
   405 => (x"87",x"c7",x"05",x"aa"),
   406 => (x"bf",x"d6",x"df",x"c2"),
   407 => (x"ca",x"87",x"cc",x"4b"),
   408 => (x"02",x"aa",x"d5",x"e9"),
   409 => (x"48",x"c0",x"87",x"c5"),
   410 => (x"c2",x"87",x"c6",x"c7"),
   411 => (x"73",x"1e",x"d0",x"d8"),
   412 => (x"87",x"df",x"f7",x"49"),
   413 => (x"98",x"70",x"86",x"c4"),
   414 => (x"c0",x"87",x"c5",x"05"),
   415 => (x"87",x"f1",x"c6",x"48"),
   416 => (x"e1",x"c0",x"1e",x"c8"),
   417 => (x"d9",x"c2",x"1e",x"cf"),
   418 => (x"d2",x"fc",x"49",x"e2"),
   419 => (x"70",x"86",x"c8",x"87"),
   420 => (x"87",x"c8",x"05",x"98"),
   421 => (x"48",x"d8",x"e0",x"c2"),
   422 => (x"87",x"da",x"78",x"c1"),
   423 => (x"e1",x"c0",x"1e",x"c8"),
   424 => (x"d9",x"c2",x"1e",x"d8"),
   425 => (x"f6",x"fb",x"49",x"c6"),
   426 => (x"70",x"86",x"c8",x"87"),
   427 => (x"c5",x"c0",x"02",x"98"),
   428 => (x"c5",x"48",x"c0",x"87"),
   429 => (x"e0",x"c2",x"87",x"fb"),
   430 => (x"49",x"bf",x"97",x"ce"),
   431 => (x"05",x"a9",x"d5",x"c1"),
   432 => (x"c2",x"87",x"cd",x"c0"),
   433 => (x"bf",x"97",x"cf",x"e0"),
   434 => (x"a9",x"ea",x"c2",x"49"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dc",x"c5",x"48",x"c0"),
   437 => (x"d0",x"d8",x"c2",x"87"),
   438 => (x"c3",x"4c",x"bf",x"97"),
   439 => (x"c0",x"02",x"ac",x"e9"),
   440 => (x"eb",x"c3",x"87",x"cc"),
   441 => (x"c5",x"c0",x"02",x"ac"),
   442 => (x"c5",x"48",x"c0",x"87"),
   443 => (x"d8",x"c2",x"87",x"c3"),
   444 => (x"49",x"bf",x"97",x"db"),
   445 => (x"cc",x"c0",x"05",x"99"),
   446 => (x"dc",x"d8",x"c2",x"87"),
   447 => (x"c2",x"49",x"bf",x"97"),
   448 => (x"c5",x"c0",x"02",x"a9"),
   449 => (x"c4",x"48",x"c0",x"87"),
   450 => (x"d8",x"c2",x"87",x"e7"),
   451 => (x"48",x"bf",x"97",x"dd"),
   452 => (x"58",x"d4",x"e0",x"c2"),
   453 => (x"e0",x"c2",x"88",x"c1"),
   454 => (x"d8",x"c2",x"58",x"d8"),
   455 => (x"49",x"bf",x"97",x"de"),
   456 => (x"d8",x"c2",x"81",x"73"),
   457 => (x"4a",x"bf",x"97",x"df"),
   458 => (x"71",x"35",x"c8",x"4d"),
   459 => (x"f0",x"e4",x"c2",x"85"),
   460 => (x"e0",x"d8",x"c2",x"5d"),
   461 => (x"c2",x"48",x"bf",x"97"),
   462 => (x"c2",x"58",x"c4",x"e5"),
   463 => (x"02",x"bf",x"d8",x"e0"),
   464 => (x"c8",x"87",x"dc",x"c2"),
   465 => (x"f4",x"e0",x"c0",x"1e"),
   466 => (x"e2",x"d9",x"c2",x"1e"),
   467 => (x"87",x"cf",x"f9",x"49"),
   468 => (x"98",x"70",x"86",x"c8"),
   469 => (x"87",x"c5",x"c0",x"02"),
   470 => (x"d4",x"c3",x"48",x"c0"),
   471 => (x"d0",x"e0",x"c2",x"87"),
   472 => (x"c4",x"48",x"4a",x"bf"),
   473 => (x"e0",x"e0",x"c2",x"30"),
   474 => (x"c0",x"e5",x"c2",x"58"),
   475 => (x"f5",x"d8",x"c2",x"5a"),
   476 => (x"c8",x"49",x"bf",x"97"),
   477 => (x"f4",x"d8",x"c2",x"31"),
   478 => (x"a1",x"4b",x"bf",x"97"),
   479 => (x"f6",x"d8",x"c2",x"49"),
   480 => (x"d0",x"4b",x"bf",x"97"),
   481 => (x"49",x"a1",x"73",x"33"),
   482 => (x"97",x"f7",x"d8",x"c2"),
   483 => (x"33",x"d8",x"4b",x"bf"),
   484 => (x"c2",x"49",x"a1",x"73"),
   485 => (x"c2",x"59",x"c8",x"e5"),
   486 => (x"91",x"bf",x"c0",x"e5"),
   487 => (x"bf",x"ec",x"e4",x"c2"),
   488 => (x"f4",x"e4",x"c2",x"81"),
   489 => (x"fd",x"d8",x"c2",x"59"),
   490 => (x"c8",x"4b",x"bf",x"97"),
   491 => (x"fc",x"d8",x"c2",x"33"),
   492 => (x"a3",x"4c",x"bf",x"97"),
   493 => (x"fe",x"d8",x"c2",x"4b"),
   494 => (x"d0",x"4c",x"bf",x"97"),
   495 => (x"4b",x"a3",x"74",x"34"),
   496 => (x"97",x"ff",x"d8",x"c2"),
   497 => (x"9c",x"cf",x"4c",x"bf"),
   498 => (x"a3",x"74",x"34",x"d8"),
   499 => (x"f8",x"e4",x"c2",x"4b"),
   500 => (x"73",x"8b",x"c2",x"5b"),
   501 => (x"f8",x"e4",x"c2",x"92"),
   502 => (x"78",x"a1",x"72",x"48"),
   503 => (x"c2",x"87",x"cb",x"c1"),
   504 => (x"bf",x"97",x"e2",x"d8"),
   505 => (x"c2",x"31",x"c8",x"49"),
   506 => (x"bf",x"97",x"e1",x"d8"),
   507 => (x"c2",x"49",x"a1",x"4a"),
   508 => (x"c5",x"59",x"e0",x"e0"),
   509 => (x"81",x"ff",x"c7",x"31"),
   510 => (x"e5",x"c2",x"29",x"c9"),
   511 => (x"d8",x"c2",x"59",x"c0"),
   512 => (x"4a",x"bf",x"97",x"e7"),
   513 => (x"d8",x"c2",x"32",x"c8"),
   514 => (x"4b",x"bf",x"97",x"e6"),
   515 => (x"e5",x"c2",x"4a",x"a2"),
   516 => (x"e5",x"c2",x"5a",x"c8"),
   517 => (x"75",x"92",x"bf",x"c0"),
   518 => (x"fc",x"e4",x"c2",x"82"),
   519 => (x"f4",x"e4",x"c2",x"5a"),
   520 => (x"c2",x"78",x"c0",x"48"),
   521 => (x"72",x"48",x"f0",x"e4"),
   522 => (x"49",x"c0",x"78",x"a1"),
   523 => (x"c1",x"87",x"f7",x"c7"),
   524 => (x"87",x"e5",x"f6",x"48"),
   525 => (x"33",x"54",x"41",x"46"),
   526 => (x"20",x"20",x"20",x"32"),
   527 => (x"54",x"41",x"46",x"00"),
   528 => (x"20",x"20",x"36",x"31"),
   529 => (x"41",x"46",x"00",x"20"),
   530 => (x"20",x"32",x"33",x"54"),
   531 => (x"46",x"00",x"20",x"20"),
   532 => (x"32",x"33",x"54",x"41"),
   533 => (x"00",x"20",x"20",x"20"),
   534 => (x"31",x"54",x"41",x"46"),
   535 => (x"20",x"20",x"20",x"36"),
   536 => (x"5b",x"5e",x"0e",x"00"),
   537 => (x"71",x"0e",x"5d",x"5c"),
   538 => (x"d8",x"e0",x"c2",x"4a"),
   539 => (x"87",x"cc",x"02",x"bf"),
   540 => (x"b7",x"c7",x"4b",x"72"),
   541 => (x"c1",x"4d",x"72",x"2b"),
   542 => (x"87",x"ca",x"9d",x"ff"),
   543 => (x"b7",x"c8",x"4b",x"72"),
   544 => (x"c3",x"4d",x"72",x"2b"),
   545 => (x"d8",x"c2",x"9d",x"ff"),
   546 => (x"e4",x"c2",x"1e",x"d0"),
   547 => (x"73",x"49",x"bf",x"ec"),
   548 => (x"fe",x"ee",x"71",x"81"),
   549 => (x"70",x"86",x"c4",x"87"),
   550 => (x"87",x"c5",x"05",x"98"),
   551 => (x"e6",x"c0",x"48",x"c0"),
   552 => (x"d8",x"e0",x"c2",x"87"),
   553 => (x"87",x"d2",x"02",x"bf"),
   554 => (x"91",x"c4",x"49",x"75"),
   555 => (x"81",x"d0",x"d8",x"c2"),
   556 => (x"ff",x"cf",x"4c",x"69"),
   557 => (x"9c",x"ff",x"ff",x"ff"),
   558 => (x"49",x"75",x"87",x"cb"),
   559 => (x"d8",x"c2",x"91",x"c2"),
   560 => (x"69",x"9f",x"81",x"d0"),
   561 => (x"f4",x"48",x"74",x"4c"),
   562 => (x"5e",x"0e",x"87",x"cf"),
   563 => (x"0e",x"5d",x"5c",x"5b"),
   564 => (x"4c",x"71",x"86",x"f4"),
   565 => (x"e5",x"c2",x"4b",x"c0"),
   566 => (x"c4",x"7e",x"bf",x"c8"),
   567 => (x"e5",x"c2",x"48",x"a6"),
   568 => (x"c8",x"78",x"bf",x"cc"),
   569 => (x"78",x"c0",x"48",x"a6"),
   570 => (x"bf",x"dc",x"e0",x"c2"),
   571 => (x"06",x"a8",x"c0",x"48"),
   572 => (x"c8",x"87",x"dd",x"c2"),
   573 => (x"99",x"cf",x"49",x"66"),
   574 => (x"c2",x"87",x"d8",x"05"),
   575 => (x"c8",x"1e",x"d0",x"d8"),
   576 => (x"c1",x"48",x"49",x"66"),
   577 => (x"58",x"a6",x"cc",x"80"),
   578 => (x"c4",x"87",x"c8",x"ed"),
   579 => (x"d0",x"d8",x"c2",x"86"),
   580 => (x"c0",x"87",x"c3",x"4b"),
   581 => (x"6b",x"97",x"83",x"e0"),
   582 => (x"c1",x"02",x"9a",x"4a"),
   583 => (x"e5",x"c3",x"87",x"e1"),
   584 => (x"da",x"c1",x"02",x"aa"),
   585 => (x"49",x"a3",x"cb",x"87"),
   586 => (x"d8",x"49",x"69",x"97"),
   587 => (x"ce",x"c1",x"05",x"99"),
   588 => (x"c0",x"1e",x"cb",x"87"),
   589 => (x"73",x"1e",x"66",x"e0"),
   590 => (x"87",x"e3",x"f1",x"49"),
   591 => (x"98",x"70",x"86",x"c8"),
   592 => (x"87",x"fb",x"c0",x"05"),
   593 => (x"c4",x"4a",x"a3",x"dc"),
   594 => (x"79",x"6a",x"49",x"a4"),
   595 => (x"c8",x"49",x"a3",x"da"),
   596 => (x"69",x"9f",x"4d",x"a4"),
   597 => (x"e0",x"c2",x"7d",x"48"),
   598 => (x"d3",x"02",x"bf",x"d8"),
   599 => (x"49",x"a3",x"d4",x"87"),
   600 => (x"c0",x"49",x"69",x"9f"),
   601 => (x"71",x"99",x"ff",x"ff"),
   602 => (x"c4",x"30",x"d0",x"48"),
   603 => (x"87",x"c2",x"58",x"a6"),
   604 => (x"48",x"6e",x"7e",x"c0"),
   605 => (x"7d",x"70",x"80",x"6d"),
   606 => (x"48",x"c1",x"7c",x"c0"),
   607 => (x"c8",x"87",x"c5",x"c1"),
   608 => (x"80",x"c1",x"48",x"66"),
   609 => (x"c2",x"58",x"a6",x"cc"),
   610 => (x"a8",x"bf",x"dc",x"e0"),
   611 => (x"87",x"e3",x"fd",x"04"),
   612 => (x"bf",x"d8",x"e0",x"c2"),
   613 => (x"87",x"ea",x"c0",x"02"),
   614 => (x"c4",x"fb",x"49",x"6e"),
   615 => (x"58",x"a6",x"c4",x"87"),
   616 => (x"ff",x"cf",x"49",x"70"),
   617 => (x"99",x"f8",x"ff",x"ff"),
   618 => (x"87",x"d6",x"02",x"a9"),
   619 => (x"89",x"c2",x"49",x"70"),
   620 => (x"bf",x"d0",x"e0",x"c2"),
   621 => (x"f0",x"e4",x"c2",x"91"),
   622 => (x"80",x"71",x"48",x"bf"),
   623 => (x"fc",x"58",x"a6",x"c8"),
   624 => (x"48",x"c0",x"87",x"e1"),
   625 => (x"d0",x"f0",x"8e",x"f4"),
   626 => (x"1e",x"73",x"1e",x"87"),
   627 => (x"49",x"6a",x"4a",x"71"),
   628 => (x"7a",x"71",x"81",x"c1"),
   629 => (x"bf",x"d4",x"e0",x"c2"),
   630 => (x"87",x"cb",x"05",x"99"),
   631 => (x"6b",x"4b",x"a2",x"c8"),
   632 => (x"87",x"fd",x"f9",x"49"),
   633 => (x"c1",x"7b",x"49",x"70"),
   634 => (x"87",x"f1",x"ef",x"48"),
   635 => (x"71",x"1e",x"73",x"1e"),
   636 => (x"f0",x"e4",x"c2",x"4b"),
   637 => (x"a3",x"c8",x"49",x"bf"),
   638 => (x"c2",x"4a",x"6a",x"4a"),
   639 => (x"d0",x"e0",x"c2",x"8a"),
   640 => (x"a1",x"72",x"92",x"bf"),
   641 => (x"d4",x"e0",x"c2",x"49"),
   642 => (x"9a",x"6b",x"4a",x"bf"),
   643 => (x"c8",x"49",x"a1",x"72"),
   644 => (x"e8",x"71",x"1e",x"66"),
   645 => (x"86",x"c4",x"87",x"fd"),
   646 => (x"c4",x"05",x"98",x"70"),
   647 => (x"c2",x"48",x"c0",x"87"),
   648 => (x"ee",x"48",x"c1",x"87"),
   649 => (x"5e",x"0e",x"87",x"f7"),
   650 => (x"71",x"0e",x"5c",x"5b"),
   651 => (x"72",x"4b",x"c0",x"4a"),
   652 => (x"e0",x"c0",x"02",x"9a"),
   653 => (x"49",x"a2",x"da",x"87"),
   654 => (x"c2",x"4b",x"69",x"9f"),
   655 => (x"02",x"bf",x"d8",x"e0"),
   656 => (x"a2",x"d4",x"87",x"cf"),
   657 => (x"49",x"69",x"9f",x"49"),
   658 => (x"ff",x"ff",x"c0",x"4c"),
   659 => (x"c2",x"34",x"d0",x"9c"),
   660 => (x"74",x"4c",x"c0",x"87"),
   661 => (x"02",x"9b",x"73",x"b3"),
   662 => (x"c2",x"4a",x"87",x"df"),
   663 => (x"d0",x"e0",x"c2",x"8a"),
   664 => (x"c2",x"92",x"49",x"bf"),
   665 => (x"48",x"bf",x"f0",x"e4"),
   666 => (x"e5",x"c2",x"80",x"72"),
   667 => (x"48",x"71",x"58",x"d0"),
   668 => (x"e0",x"c2",x"30",x"c4"),
   669 => (x"e9",x"c0",x"58",x"e0"),
   670 => (x"f4",x"e4",x"c2",x"87"),
   671 => (x"e5",x"c2",x"4b",x"bf"),
   672 => (x"e4",x"c2",x"48",x"cc"),
   673 => (x"c2",x"78",x"bf",x"f8"),
   674 => (x"02",x"bf",x"d8",x"e0"),
   675 => (x"e0",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"d0"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"fc",x"e4"),
   679 => (x"e0",x"c2",x"31",x"c4"),
   680 => (x"e5",x"c2",x"59",x"e0"),
   681 => (x"f2",x"ec",x"5b",x"cc"),
   682 => (x"5b",x"5e",x"0e",x"87"),
   683 => (x"f4",x"0e",x"5d",x"5c"),
   684 => (x"9a",x"4a",x"71",x"86"),
   685 => (x"c2",x"87",x"de",x"02"),
   686 => (x"c0",x"48",x"cc",x"d8"),
   687 => (x"c4",x"d8",x"c2",x"78"),
   688 => (x"cc",x"e5",x"c2",x"48"),
   689 => (x"d8",x"c2",x"78",x"bf"),
   690 => (x"e5",x"c2",x"48",x"c8"),
   691 => (x"c0",x"78",x"bf",x"c8"),
   692 => (x"c0",x"48",x"ff",x"f1"),
   693 => (x"dc",x"e0",x"c2",x"78"),
   694 => (x"d8",x"c2",x"49",x"bf"),
   695 => (x"71",x"4a",x"bf",x"cc"),
   696 => (x"cb",x"c4",x"03",x"aa"),
   697 => (x"cf",x"49",x"72",x"87"),
   698 => (x"e0",x"c0",x"05",x"99"),
   699 => (x"d0",x"d8",x"c2",x"87"),
   700 => (x"c4",x"d8",x"c2",x"1e"),
   701 => (x"d8",x"c2",x"49",x"bf"),
   702 => (x"a1",x"c1",x"48",x"c4"),
   703 => (x"d2",x"e5",x"71",x"78"),
   704 => (x"c0",x"86",x"c4",x"87"),
   705 => (x"c2",x"48",x"fb",x"f1"),
   706 => (x"cc",x"78",x"d0",x"d8"),
   707 => (x"fb",x"f1",x"c0",x"87"),
   708 => (x"e0",x"c0",x"48",x"bf"),
   709 => (x"ff",x"f1",x"c0",x"80"),
   710 => (x"cc",x"d8",x"c2",x"58"),
   711 => (x"80",x"c1",x"48",x"bf"),
   712 => (x"58",x"d0",x"d8",x"c2"),
   713 => (x"00",x"0c",x"7b",x"27"),
   714 => (x"bf",x"97",x"bf",x"00"),
   715 => (x"c2",x"02",x"9c",x"4c"),
   716 => (x"e5",x"c3",x"87",x"ee"),
   717 => (x"e7",x"c2",x"02",x"ac"),
   718 => (x"fb",x"f1",x"c0",x"87"),
   719 => (x"a3",x"cb",x"4b",x"bf"),
   720 => (x"cf",x"4d",x"11",x"49"),
   721 => (x"d6",x"c1",x"05",x"ad"),
   722 => (x"df",x"49",x"74",x"87"),
   723 => (x"cd",x"89",x"c1",x"99"),
   724 => (x"e0",x"e0",x"c2",x"91"),
   725 => (x"4a",x"a3",x"c1",x"81"),
   726 => (x"a3",x"c3",x"51",x"12"),
   727 => (x"c5",x"51",x"12",x"4a"),
   728 => (x"51",x"12",x"4a",x"a3"),
   729 => (x"12",x"4a",x"a3",x"c7"),
   730 => (x"4a",x"a3",x"c9",x"51"),
   731 => (x"a3",x"ce",x"51",x"12"),
   732 => (x"d0",x"51",x"12",x"4a"),
   733 => (x"51",x"12",x"4a",x"a3"),
   734 => (x"12",x"4a",x"a3",x"d2"),
   735 => (x"4a",x"a3",x"d4",x"51"),
   736 => (x"a3",x"d6",x"51",x"12"),
   737 => (x"d8",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"dc"),
   740 => (x"4a",x"a3",x"de",x"51"),
   741 => (x"f1",x"c0",x"51",x"12"),
   742 => (x"78",x"c1",x"48",x"ff"),
   743 => (x"75",x"87",x"c1",x"c1"),
   744 => (x"05",x"99",x"c8",x"49"),
   745 => (x"75",x"87",x"f3",x"c0"),
   746 => (x"05",x"99",x"d0",x"49"),
   747 => (x"66",x"dc",x"87",x"d0"),
   748 => (x"87",x"ca",x"c0",x"02"),
   749 => (x"66",x"dc",x"49",x"73"),
   750 => (x"02",x"98",x"70",x"0f"),
   751 => (x"f1",x"c0",x"87",x"dc"),
   752 => (x"c0",x"05",x"bf",x"ff"),
   753 => (x"e0",x"c2",x"87",x"c6"),
   754 => (x"50",x"c0",x"48",x"e0"),
   755 => (x"48",x"ff",x"f1",x"c0"),
   756 => (x"f1",x"c0",x"78",x"c0"),
   757 => (x"c2",x"48",x"bf",x"fb"),
   758 => (x"f1",x"c0",x"87",x"dc"),
   759 => (x"78",x"c0",x"48",x"ff"),
   760 => (x"bf",x"dc",x"e0",x"c2"),
   761 => (x"cc",x"d8",x"c2",x"49"),
   762 => (x"aa",x"71",x"4a",x"bf"),
   763 => (x"87",x"f5",x"fb",x"04"),
   764 => (x"bf",x"cc",x"e5",x"c2"),
   765 => (x"87",x"c8",x"c0",x"05"),
   766 => (x"bf",x"d8",x"e0",x"c2"),
   767 => (x"87",x"f4",x"c1",x"02"),
   768 => (x"bf",x"c8",x"d8",x"c2"),
   769 => (x"87",x"d9",x"f1",x"49"),
   770 => (x"58",x"cc",x"d8",x"c2"),
   771 => (x"e0",x"c2",x"7e",x"70"),
   772 => (x"c0",x"02",x"bf",x"d8"),
   773 => (x"49",x"6e",x"87",x"dd"),
   774 => (x"ff",x"ff",x"ff",x"cf"),
   775 => (x"02",x"a9",x"99",x"f8"),
   776 => (x"c4",x"87",x"c8",x"c0"),
   777 => (x"78",x"c0",x"48",x"a6"),
   778 => (x"c4",x"87",x"e6",x"c0"),
   779 => (x"78",x"c1",x"48",x"a6"),
   780 => (x"6e",x"87",x"de",x"c0"),
   781 => (x"f8",x"ff",x"cf",x"49"),
   782 => (x"c0",x"02",x"a9",x"99"),
   783 => (x"a6",x"c8",x"87",x"c8"),
   784 => (x"c0",x"78",x"c0",x"48"),
   785 => (x"a6",x"c8",x"87",x"c5"),
   786 => (x"c4",x"78",x"c1",x"48"),
   787 => (x"66",x"c8",x"48",x"a6"),
   788 => (x"05",x"66",x"c4",x"78"),
   789 => (x"6e",x"87",x"dd",x"c0"),
   790 => (x"c2",x"89",x"c2",x"49"),
   791 => (x"91",x"bf",x"d0",x"e0"),
   792 => (x"bf",x"f0",x"e4",x"c2"),
   793 => (x"c2",x"80",x"71",x"48"),
   794 => (x"c2",x"58",x"c8",x"d8"),
   795 => (x"c0",x"48",x"cc",x"d8"),
   796 => (x"87",x"e1",x"f9",x"78"),
   797 => (x"8e",x"f4",x"48",x"c0"),
   798 => (x"00",x"87",x"de",x"e5"),
   799 => (x"00",x"00",x"00",x"00"),
   800 => (x"1e",x"00",x"00",x"00"),
   801 => (x"c3",x"48",x"d4",x"ff"),
   802 => (x"49",x"68",x"78",x"ff"),
   803 => (x"87",x"c6",x"02",x"99"),
   804 => (x"05",x"a9",x"fb",x"c0"),
   805 => (x"48",x"71",x"87",x"ee"),
   806 => (x"5e",x"0e",x"4f",x"26"),
   807 => (x"71",x"0e",x"5c",x"5b"),
   808 => (x"ff",x"4b",x"c0",x"4a"),
   809 => (x"ff",x"c3",x"48",x"d4"),
   810 => (x"99",x"49",x"68",x"78"),
   811 => (x"87",x"c1",x"c1",x"02"),
   812 => (x"02",x"a9",x"ec",x"c0"),
   813 => (x"c0",x"87",x"fa",x"c0"),
   814 => (x"c0",x"02",x"a9",x"fb"),
   815 => (x"66",x"cc",x"87",x"f3"),
   816 => (x"cc",x"03",x"ab",x"b7"),
   817 => (x"02",x"66",x"d0",x"87"),
   818 => (x"09",x"72",x"87",x"c7"),
   819 => (x"c1",x"09",x"79",x"97"),
   820 => (x"02",x"99",x"71",x"82"),
   821 => (x"83",x"c1",x"87",x"c2"),
   822 => (x"c3",x"48",x"d4",x"ff"),
   823 => (x"49",x"68",x"78",x"ff"),
   824 => (x"87",x"cd",x"02",x"99"),
   825 => (x"02",x"a9",x"ec",x"c0"),
   826 => (x"fb",x"c0",x"87",x"c7"),
   827 => (x"cd",x"ff",x"05",x"a9"),
   828 => (x"02",x"66",x"d0",x"87"),
   829 => (x"97",x"c0",x"87",x"c3"),
   830 => (x"a9",x"fb",x"c0",x"7a"),
   831 => (x"73",x"87",x"c7",x"05"),
   832 => (x"8c",x"0c",x"c0",x"4c"),
   833 => (x"4c",x"73",x"87",x"c2"),
   834 => (x"87",x"c2",x"48",x"74"),
   835 => (x"4c",x"26",x"4d",x"26"),
   836 => (x"4f",x"26",x"4b",x"26"),
   837 => (x"48",x"d4",x"ff",x"1e"),
   838 => (x"68",x"78",x"ff",x"c3"),
   839 => (x"b7",x"f0",x"c0",x"49"),
   840 => (x"87",x"ca",x"04",x"a9"),
   841 => (x"a9",x"b7",x"f9",x"c0"),
   842 => (x"c0",x"87",x"c3",x"01"),
   843 => (x"c1",x"c1",x"89",x"f0"),
   844 => (x"ca",x"04",x"a9",x"b7"),
   845 => (x"b7",x"c6",x"c1",x"87"),
   846 => (x"87",x"c3",x"01",x"a9"),
   847 => (x"71",x"89",x"f7",x"c0"),
   848 => (x"0e",x"4f",x"26",x"48"),
   849 => (x"5d",x"5c",x"5b",x"5e"),
   850 => (x"71",x"86",x"f4",x"0e"),
   851 => (x"4b",x"d4",x"ff",x"4c"),
   852 => (x"c3",x"7e",x"4d",x"c0"),
   853 => (x"d0",x"ff",x"7b",x"ff"),
   854 => (x"c0",x"c8",x"48",x"bf"),
   855 => (x"a6",x"c8",x"98",x"c0"),
   856 => (x"02",x"98",x"70",x"58"),
   857 => (x"d0",x"ff",x"87",x"d0"),
   858 => (x"c0",x"c8",x"48",x"bf"),
   859 => (x"a6",x"c8",x"98",x"c0"),
   860 => (x"05",x"98",x"70",x"58"),
   861 => (x"d0",x"ff",x"87",x"f0"),
   862 => (x"78",x"e1",x"c0",x"48"),
   863 => (x"c2",x"fc",x"7b",x"d4"),
   864 => (x"99",x"49",x"70",x"87"),
   865 => (x"87",x"c7",x"c1",x"02"),
   866 => (x"c8",x"7b",x"ff",x"c3"),
   867 => (x"78",x"6b",x"48",x"a6"),
   868 => (x"c0",x"48",x"66",x"c8"),
   869 => (x"c8",x"02",x"a8",x"fb"),
   870 => (x"e8",x"e5",x"c2",x"87"),
   871 => (x"ee",x"c0",x"02",x"bf"),
   872 => (x"71",x"4d",x"c1",x"87"),
   873 => (x"e6",x"c0",x"02",x"99"),
   874 => (x"a9",x"fb",x"c0",x"87"),
   875 => (x"fb",x"87",x"c3",x"02"),
   876 => (x"ff",x"c3",x"87",x"d1"),
   877 => (x"c1",x"49",x"6b",x"7b"),
   878 => (x"cc",x"05",x"a9",x"c6"),
   879 => (x"7b",x"ff",x"c3",x"87"),
   880 => (x"48",x"a6",x"c8",x"7b"),
   881 => (x"49",x"c0",x"78",x"6b"),
   882 => (x"05",x"99",x"71",x"4d"),
   883 => (x"75",x"87",x"da",x"ff"),
   884 => (x"de",x"c1",x"05",x"9d"),
   885 => (x"7b",x"ff",x"c3",x"87"),
   886 => (x"ff",x"c3",x"4a",x"6b"),
   887 => (x"48",x"a6",x"c4",x"7b"),
   888 => (x"48",x"6e",x"78",x"6b"),
   889 => (x"a6",x"c4",x"80",x"c1"),
   890 => (x"49",x"a4",x"c8",x"58"),
   891 => (x"c8",x"49",x"69",x"97"),
   892 => (x"da",x"05",x"a9",x"66"),
   893 => (x"49",x"a4",x"c9",x"87"),
   894 => (x"aa",x"49",x"69",x"97"),
   895 => (x"ca",x"87",x"d0",x"05"),
   896 => (x"69",x"97",x"49",x"a4"),
   897 => (x"a9",x"66",x"c4",x"49"),
   898 => (x"c1",x"87",x"c4",x"05"),
   899 => (x"c8",x"87",x"d6",x"4d"),
   900 => (x"ec",x"c0",x"48",x"66"),
   901 => (x"87",x"c9",x"02",x"a8"),
   902 => (x"c0",x"48",x"66",x"c8"),
   903 => (x"c4",x"05",x"a8",x"fb"),
   904 => (x"c1",x"7e",x"c0",x"87"),
   905 => (x"7b",x"ff",x"c3",x"4d"),
   906 => (x"6b",x"48",x"a6",x"c8"),
   907 => (x"02",x"9d",x"75",x"78"),
   908 => (x"ff",x"87",x"e2",x"fe"),
   909 => (x"c8",x"48",x"bf",x"d0"),
   910 => (x"c8",x"98",x"c0",x"c0"),
   911 => (x"98",x"70",x"58",x"a6"),
   912 => (x"ff",x"87",x"d0",x"02"),
   913 => (x"c8",x"48",x"bf",x"d0"),
   914 => (x"c8",x"98",x"c0",x"c0"),
   915 => (x"98",x"70",x"58",x"a6"),
   916 => (x"ff",x"87",x"f0",x"05"),
   917 => (x"e0",x"c0",x"48",x"d0"),
   918 => (x"f4",x"48",x"6e",x"78"),
   919 => (x"87",x"ec",x"fa",x"8e"),
   920 => (x"5c",x"5b",x"5e",x"0e"),
   921 => (x"86",x"f4",x"0e",x"5d"),
   922 => (x"ff",x"59",x"a6",x"c4"),
   923 => (x"c0",x"c8",x"4c",x"d0"),
   924 => (x"1e",x"6e",x"4b",x"c0"),
   925 => (x"49",x"ec",x"e5",x"c2"),
   926 => (x"c4",x"87",x"cf",x"e9"),
   927 => (x"02",x"98",x"70",x"86"),
   928 => (x"c2",x"87",x"f7",x"c5"),
   929 => (x"4d",x"bf",x"f0",x"e5"),
   930 => (x"f6",x"fa",x"49",x"6e"),
   931 => (x"58",x"a6",x"c8",x"87"),
   932 => (x"98",x"73",x"48",x"6c"),
   933 => (x"70",x"58",x"a6",x"cc"),
   934 => (x"87",x"cc",x"02",x"98"),
   935 => (x"98",x"73",x"48",x"6c"),
   936 => (x"70",x"58",x"a6",x"c4"),
   937 => (x"87",x"f4",x"05",x"98"),
   938 => (x"d4",x"ff",x"7c",x"c5"),
   939 => (x"78",x"d5",x"c1",x"48"),
   940 => (x"bf",x"e8",x"e5",x"c2"),
   941 => (x"c4",x"81",x"c1",x"49"),
   942 => (x"8a",x"c1",x"4a",x"66"),
   943 => (x"48",x"72",x"32",x"c6"),
   944 => (x"d4",x"ff",x"b0",x"71"),
   945 => (x"48",x"6c",x"78",x"08"),
   946 => (x"a6",x"c4",x"98",x"73"),
   947 => (x"02",x"98",x"70",x"58"),
   948 => (x"48",x"6c",x"87",x"cc"),
   949 => (x"a6",x"c4",x"98",x"73"),
   950 => (x"05",x"98",x"70",x"58"),
   951 => (x"7c",x"c4",x"87",x"f4"),
   952 => (x"c3",x"48",x"d4",x"ff"),
   953 => (x"48",x"6c",x"78",x"ff"),
   954 => (x"a6",x"c4",x"98",x"73"),
   955 => (x"02",x"98",x"70",x"58"),
   956 => (x"48",x"6c",x"87",x"cc"),
   957 => (x"a6",x"c4",x"98",x"73"),
   958 => (x"05",x"98",x"70",x"58"),
   959 => (x"7c",x"c5",x"87",x"f4"),
   960 => (x"c1",x"48",x"d4",x"ff"),
   961 => (x"78",x"c1",x"78",x"d3"),
   962 => (x"98",x"73",x"48",x"6c"),
   963 => (x"70",x"58",x"a6",x"c4"),
   964 => (x"87",x"cc",x"02",x"98"),
   965 => (x"98",x"73",x"48",x"6c"),
   966 => (x"70",x"58",x"a6",x"c4"),
   967 => (x"87",x"f4",x"05",x"98"),
   968 => (x"9d",x"75",x"7c",x"c4"),
   969 => (x"87",x"d0",x"c2",x"02"),
   970 => (x"7e",x"d0",x"d8",x"c2"),
   971 => (x"ec",x"e5",x"c2",x"1e"),
   972 => (x"87",x"f8",x"ea",x"49"),
   973 => (x"98",x"70",x"86",x"c4"),
   974 => (x"c0",x"87",x"c5",x"05"),
   975 => (x"87",x"fc",x"c2",x"48"),
   976 => (x"ad",x"b7",x"c0",x"c8"),
   977 => (x"4a",x"87",x"c4",x"04"),
   978 => (x"75",x"87",x"c4",x"8d"),
   979 => (x"6c",x"4d",x"c0",x"4a"),
   980 => (x"c8",x"98",x"73",x"48"),
   981 => (x"98",x"70",x"58",x"a6"),
   982 => (x"6c",x"87",x"cc",x"02"),
   983 => (x"c8",x"98",x"73",x"48"),
   984 => (x"98",x"70",x"58",x"a6"),
   985 => (x"cd",x"87",x"f4",x"05"),
   986 => (x"48",x"d4",x"ff",x"7c"),
   987 => (x"72",x"78",x"d4",x"c1"),
   988 => (x"71",x"8a",x"c1",x"49"),
   989 => (x"87",x"d9",x"02",x"99"),
   990 => (x"48",x"bf",x"97",x"6e"),
   991 => (x"78",x"08",x"d4",x"ff"),
   992 => (x"80",x"c1",x"48",x"6e"),
   993 => (x"72",x"58",x"a6",x"c4"),
   994 => (x"71",x"8a",x"c1",x"49"),
   995 => (x"e7",x"ff",x"05",x"99"),
   996 => (x"73",x"48",x"6c",x"87"),
   997 => (x"58",x"a6",x"c4",x"98"),
   998 => (x"cc",x"02",x"98",x"70"),
   999 => (x"73",x"48",x"6c",x"87"),
  1000 => (x"58",x"a6",x"c4",x"98"),
  1001 => (x"f4",x"05",x"98",x"70"),
  1002 => (x"c2",x"7c",x"c4",x"87"),
  1003 => (x"e8",x"49",x"ec",x"e5"),
  1004 => (x"9d",x"75",x"87",x"d7"),
  1005 => (x"87",x"f0",x"fd",x"05"),
  1006 => (x"98",x"73",x"48",x"6c"),
  1007 => (x"70",x"58",x"a6",x"c4"),
  1008 => (x"87",x"cd",x"02",x"98"),
  1009 => (x"98",x"73",x"48",x"6c"),
  1010 => (x"70",x"58",x"a6",x"c4"),
  1011 => (x"f3",x"ff",x"05",x"98"),
  1012 => (x"ff",x"7c",x"c5",x"87"),
  1013 => (x"d3",x"c1",x"48",x"d4"),
  1014 => (x"6c",x"78",x"c0",x"78"),
  1015 => (x"c4",x"98",x"73",x"48"),
  1016 => (x"98",x"70",x"58",x"a6"),
  1017 => (x"6c",x"87",x"cd",x"02"),
  1018 => (x"c4",x"98",x"73",x"48"),
  1019 => (x"98",x"70",x"58",x"a6"),
  1020 => (x"87",x"f3",x"ff",x"05"),
  1021 => (x"48",x"c1",x"7c",x"c4"),
  1022 => (x"48",x"c0",x"87",x"c2"),
  1023 => (x"cb",x"f4",x"8e",x"f4"),
  1024 => (x"5b",x"5e",x"0e",x"87"),
  1025 => (x"1e",x"0e",x"5d",x"5c"),
  1026 => (x"4c",x"c0",x"4b",x"71"),
  1027 => (x"04",x"ab",x"b7",x"4d"),
  1028 => (x"c0",x"87",x"e9",x"c0"),
  1029 => (x"75",x"1e",x"c3",x"f5"),
  1030 => (x"87",x"c4",x"02",x"9d"),
  1031 => (x"87",x"c2",x"4a",x"c0"),
  1032 => (x"49",x"72",x"4a",x"c1"),
  1033 => (x"c4",x"87",x"c2",x"ea"),
  1034 => (x"c1",x"58",x"a6",x"86"),
  1035 => (x"c2",x"05",x"6e",x"84"),
  1036 => (x"c1",x"4c",x"73",x"87"),
  1037 => (x"ac",x"b7",x"73",x"85"),
  1038 => (x"87",x"d7",x"ff",x"06"),
  1039 => (x"f3",x"26",x"48",x"6e"),
  1040 => (x"5e",x"0e",x"87",x"ca"),
  1041 => (x"0e",x"5d",x"5c",x"5b"),
  1042 => (x"49",x"4c",x"71",x"1e"),
  1043 => (x"bf",x"fc",x"e5",x"c2"),
  1044 => (x"87",x"ed",x"fe",x"81"),
  1045 => (x"02",x"9d",x"4d",x"70"),
  1046 => (x"c2",x"87",x"fc",x"c0"),
  1047 => (x"75",x"4b",x"e0",x"e0"),
  1048 => (x"ff",x"49",x"cb",x"4a"),
  1049 => (x"74",x"87",x"c9",x"c1"),
  1050 => (x"c2",x"91",x"de",x"49"),
  1051 => (x"71",x"48",x"d0",x"e6"),
  1052 => (x"58",x"a6",x"c4",x"80"),
  1053 => (x"48",x"e7",x"c2",x"c1"),
  1054 => (x"a1",x"c8",x"49",x"6e"),
  1055 => (x"71",x"41",x"20",x"4a"),
  1056 => (x"87",x"f9",x"05",x"aa"),
  1057 => (x"51",x"10",x"51",x"10"),
  1058 => (x"49",x"74",x"51",x"10"),
  1059 => (x"87",x"ee",x"c5",x"c1"),
  1060 => (x"49",x"e0",x"e0",x"c2"),
  1061 => (x"c1",x"87",x"c9",x"f7"),
  1062 => (x"c1",x"49",x"e0",x"e4"),
  1063 => (x"c1",x"87",x"f6",x"c7"),
  1064 => (x"26",x"87",x"d2",x"c8"),
  1065 => (x"4c",x"87",x"e5",x"f1"),
  1066 => (x"69",x"64",x"61",x"6f"),
  1067 => (x"2e",x"2e",x"67",x"6e"),
  1068 => (x"20",x"80",x"00",x"2e"),
  1069 => (x"6b",x"63",x"61",x"42"),
  1070 => (x"61",x"6f",x"4c",x"00"),
  1071 => (x"2e",x"2a",x"20",x"64"),
  1072 => (x"20",x"3a",x"00",x"20"),
  1073 => (x"42",x"20",x"80",x"00"),
  1074 => (x"00",x"6b",x"63",x"61"),
  1075 => (x"78",x"45",x"20",x"80"),
  1076 => (x"53",x"00",x"74",x"69"),
  1077 => (x"6e",x"49",x"20",x"44"),
  1078 => (x"2e",x"2e",x"74",x"69"),
  1079 => (x"00",x"4b",x"4f",x"00"),
  1080 => (x"54",x"4f",x"4f",x"42"),
  1081 => (x"20",x"20",x"20",x"20"),
  1082 => (x"00",x"4d",x"4f",x"52"),
  1083 => (x"71",x"1e",x"73",x"1e"),
  1084 => (x"e5",x"c2",x"49",x"4b"),
  1085 => (x"fc",x"81",x"bf",x"fc"),
  1086 => (x"4a",x"70",x"87",x"c7"),
  1087 => (x"87",x"c4",x"02",x"9a"),
  1088 => (x"87",x"e2",x"e4",x"49"),
  1089 => (x"48",x"fc",x"e5",x"c2"),
  1090 => (x"49",x"73",x"78",x"c0"),
  1091 => (x"ef",x"87",x"e9",x"c1"),
  1092 => (x"73",x"1e",x"87",x"fe"),
  1093 => (x"c4",x"4b",x"71",x"1e"),
  1094 => (x"c1",x"02",x"4a",x"a3"),
  1095 => (x"8a",x"c1",x"87",x"c8"),
  1096 => (x"8a",x"87",x"dc",x"02"),
  1097 => (x"87",x"f1",x"c0",x"02"),
  1098 => (x"c4",x"c1",x"05",x"8a"),
  1099 => (x"fc",x"e5",x"c2",x"87"),
  1100 => (x"fc",x"c0",x"02",x"bf"),
  1101 => (x"88",x"c1",x"48",x"87"),
  1102 => (x"58",x"c0",x"e6",x"c2"),
  1103 => (x"c2",x"87",x"f2",x"c0"),
  1104 => (x"49",x"bf",x"fc",x"e5"),
  1105 => (x"e6",x"c2",x"89",x"d0"),
  1106 => (x"b7",x"c0",x"59",x"c0"),
  1107 => (x"e0",x"c0",x"03",x"a9"),
  1108 => (x"fc",x"e5",x"c2",x"87"),
  1109 => (x"d8",x"78",x"c0",x"48"),
  1110 => (x"fc",x"e5",x"c2",x"87"),
  1111 => (x"80",x"c1",x"48",x"bf"),
  1112 => (x"58",x"c0",x"e6",x"c2"),
  1113 => (x"e5",x"c2",x"87",x"cb"),
  1114 => (x"d0",x"48",x"bf",x"fc"),
  1115 => (x"c0",x"e6",x"c2",x"80"),
  1116 => (x"c3",x"49",x"73",x"58"),
  1117 => (x"87",x"d8",x"ee",x"87"),
  1118 => (x"5c",x"5b",x"5e",x"0e"),
  1119 => (x"86",x"f0",x"0e",x"5d"),
  1120 => (x"c2",x"59",x"a6",x"d0"),
  1121 => (x"c0",x"4d",x"d0",x"d8"),
  1122 => (x"48",x"a6",x"c4",x"4c"),
  1123 => (x"e5",x"c2",x"78",x"c0"),
  1124 => (x"c0",x"48",x"bf",x"fc"),
  1125 => (x"c1",x"06",x"a8",x"b7"),
  1126 => (x"d8",x"c2",x"87",x"c1"),
  1127 => (x"02",x"98",x"48",x"d0"),
  1128 => (x"c0",x"87",x"f8",x"c0"),
  1129 => (x"c8",x"1e",x"c3",x"f5"),
  1130 => (x"87",x"c7",x"02",x"66"),
  1131 => (x"c0",x"48",x"a6",x"c4"),
  1132 => (x"c4",x"87",x"c5",x"78"),
  1133 => (x"78",x"c1",x"48",x"a6"),
  1134 => (x"e3",x"49",x"66",x"c4"),
  1135 => (x"86",x"c4",x"87",x"eb"),
  1136 => (x"84",x"c1",x"4d",x"70"),
  1137 => (x"c1",x"48",x"66",x"c4"),
  1138 => (x"58",x"a6",x"c8",x"80"),
  1139 => (x"bf",x"fc",x"e5",x"c2"),
  1140 => (x"c6",x"03",x"ac",x"b7"),
  1141 => (x"05",x"9d",x"75",x"87"),
  1142 => (x"c0",x"87",x"c8",x"ff"),
  1143 => (x"02",x"9d",x"75",x"4c"),
  1144 => (x"c0",x"87",x"e3",x"c3"),
  1145 => (x"c8",x"1e",x"c3",x"f5"),
  1146 => (x"87",x"c7",x"02",x"66"),
  1147 => (x"c0",x"48",x"a6",x"cc"),
  1148 => (x"cc",x"87",x"c5",x"78"),
  1149 => (x"78",x"c1",x"48",x"a6"),
  1150 => (x"e2",x"49",x"66",x"cc"),
  1151 => (x"86",x"c4",x"87",x"eb"),
  1152 => (x"02",x"6e",x"58",x"a6"),
  1153 => (x"49",x"87",x"eb",x"c2"),
  1154 => (x"69",x"97",x"81",x"cb"),
  1155 => (x"02",x"99",x"d0",x"49"),
  1156 => (x"c1",x"87",x"d9",x"c1"),
  1157 => (x"74",x"4b",x"ec",x"c3"),
  1158 => (x"c1",x"91",x"cc",x"49"),
  1159 => (x"c8",x"81",x"e0",x"e4"),
  1160 => (x"7a",x"73",x"4a",x"a1"),
  1161 => (x"ff",x"c3",x"81",x"c1"),
  1162 => (x"de",x"49",x"74",x"51"),
  1163 => (x"d0",x"e6",x"c2",x"91"),
  1164 => (x"c2",x"85",x"71",x"4d"),
  1165 => (x"c1",x"7d",x"97",x"c1"),
  1166 => (x"e0",x"c0",x"49",x"a5"),
  1167 => (x"e0",x"e0",x"c2",x"51"),
  1168 => (x"d2",x"02",x"bf",x"97"),
  1169 => (x"c2",x"84",x"c1",x"87"),
  1170 => (x"e0",x"c2",x"4b",x"a5"),
  1171 => (x"49",x"db",x"4a",x"e0"),
  1172 => (x"87",x"dc",x"f9",x"fe"),
  1173 => (x"cd",x"87",x"db",x"c1"),
  1174 => (x"51",x"c0",x"49",x"a5"),
  1175 => (x"a5",x"c2",x"84",x"c1"),
  1176 => (x"cb",x"4a",x"6e",x"4b"),
  1177 => (x"c7",x"f9",x"fe",x"49"),
  1178 => (x"87",x"c6",x"c1",x"87"),
  1179 => (x"91",x"cc",x"49",x"74"),
  1180 => (x"81",x"e0",x"e4",x"c1"),
  1181 => (x"c1",x"c1",x"81",x"c8"),
  1182 => (x"e0",x"c2",x"79",x"c2"),
  1183 => (x"02",x"bf",x"97",x"e0"),
  1184 => (x"49",x"74",x"87",x"d8"),
  1185 => (x"84",x"c1",x"91",x"de"),
  1186 => (x"4b",x"d0",x"e6",x"c2"),
  1187 => (x"e0",x"c2",x"83",x"71"),
  1188 => (x"49",x"dd",x"4a",x"e0"),
  1189 => (x"87",x"d8",x"f8",x"fe"),
  1190 => (x"4b",x"74",x"87",x"d8"),
  1191 => (x"e6",x"c2",x"93",x"de"),
  1192 => (x"a3",x"cb",x"83",x"d0"),
  1193 => (x"c1",x"51",x"c0",x"49"),
  1194 => (x"4a",x"6e",x"73",x"84"),
  1195 => (x"f7",x"fe",x"49",x"cb"),
  1196 => (x"66",x"c4",x"87",x"fe"),
  1197 => (x"c8",x"80",x"c1",x"48"),
  1198 => (x"b7",x"c7",x"58",x"a6"),
  1199 => (x"c5",x"c0",x"03",x"ac"),
  1200 => (x"fc",x"05",x"6e",x"87"),
  1201 => (x"b7",x"c7",x"87",x"dd"),
  1202 => (x"d3",x"c0",x"03",x"ac"),
  1203 => (x"de",x"49",x"74",x"87"),
  1204 => (x"d0",x"e6",x"c2",x"91"),
  1205 => (x"c1",x"51",x"c0",x"81"),
  1206 => (x"ac",x"b7",x"c7",x"84"),
  1207 => (x"87",x"ed",x"ff",x"04"),
  1208 => (x"48",x"f5",x"e5",x"c1"),
  1209 => (x"e5",x"c1",x"50",x"c0"),
  1210 => (x"50",x"c2",x"48",x"f4"),
  1211 => (x"48",x"fc",x"e5",x"c1"),
  1212 => (x"78",x"de",x"cc",x"c1"),
  1213 => (x"48",x"f8",x"e5",x"c1"),
  1214 => (x"78",x"f2",x"c2",x"c1"),
  1215 => (x"48",x"c8",x"e6",x"c1"),
  1216 => (x"78",x"d2",x"c4",x"c1"),
  1217 => (x"c0",x"49",x"66",x"cc"),
  1218 => (x"f0",x"87",x"f3",x"fb"),
  1219 => (x"87",x"fc",x"e7",x"8e"),
  1220 => (x"c2",x"4a",x"71",x"1e"),
  1221 => (x"72",x"5a",x"ec",x"e5"),
  1222 => (x"87",x"dc",x"f9",x"49"),
  1223 => (x"71",x"1e",x"4f",x"26"),
  1224 => (x"91",x"cc",x"49",x"4a"),
  1225 => (x"81",x"e0",x"e4",x"c1"),
  1226 => (x"48",x"11",x"81",x"c1"),
  1227 => (x"58",x"e8",x"e5",x"c2"),
  1228 => (x"49",x"a2",x"f0",x"c0"),
  1229 => (x"87",x"c8",x"f6",x"fe"),
  1230 => (x"dd",x"d5",x"49",x"c0"),
  1231 => (x"0e",x"4f",x"26",x"87"),
  1232 => (x"5d",x"5c",x"5b",x"5e"),
  1233 => (x"71",x"86",x"f0",x"0e"),
  1234 => (x"91",x"cc",x"49",x"4c"),
  1235 => (x"81",x"e0",x"e4",x"c1"),
  1236 => (x"c4",x"7e",x"a1",x"c3"),
  1237 => (x"e5",x"c2",x"48",x"a6"),
  1238 => (x"6e",x"78",x"bf",x"e0"),
  1239 => (x"c4",x"4a",x"bf",x"97"),
  1240 => (x"2b",x"72",x"4b",x"66"),
  1241 => (x"12",x"4a",x"a1",x"c1"),
  1242 => (x"58",x"a6",x"cc",x"48"),
  1243 => (x"83",x"c1",x"9b",x"70"),
  1244 => (x"69",x"97",x"81",x"c2"),
  1245 => (x"04",x"ab",x"b7",x"49"),
  1246 => (x"4b",x"c0",x"87",x"c2"),
  1247 => (x"4a",x"bf",x"97",x"6e"),
  1248 => (x"72",x"49",x"66",x"c8"),
  1249 => (x"c4",x"b9",x"ff",x"31"),
  1250 => (x"4d",x"73",x"99",x"66"),
  1251 => (x"b5",x"71",x"35",x"72"),
  1252 => (x"5d",x"e4",x"e5",x"c2"),
  1253 => (x"c3",x"48",x"d4",x"ff"),
  1254 => (x"d0",x"ff",x"78",x"ff"),
  1255 => (x"c0",x"c8",x"48",x"bf"),
  1256 => (x"a6",x"d0",x"98",x"c0"),
  1257 => (x"02",x"98",x"70",x"58"),
  1258 => (x"d0",x"ff",x"87",x"d0"),
  1259 => (x"c0",x"c8",x"48",x"bf"),
  1260 => (x"a6",x"c4",x"98",x"c0"),
  1261 => (x"05",x"98",x"70",x"58"),
  1262 => (x"d0",x"ff",x"87",x"f0"),
  1263 => (x"78",x"e1",x"c0",x"48"),
  1264 => (x"de",x"48",x"d4",x"ff"),
  1265 => (x"7d",x"0d",x"70",x"78"),
  1266 => (x"c8",x"48",x"75",x"0d"),
  1267 => (x"d4",x"ff",x"28",x"b7"),
  1268 => (x"48",x"75",x"78",x"08"),
  1269 => (x"ff",x"28",x"b7",x"d0"),
  1270 => (x"75",x"78",x"08",x"d4"),
  1271 => (x"28",x"b7",x"d8",x"48"),
  1272 => (x"78",x"08",x"d4",x"ff"),
  1273 => (x"48",x"bf",x"d0",x"ff"),
  1274 => (x"98",x"c0",x"c0",x"c8"),
  1275 => (x"70",x"58",x"a6",x"c4"),
  1276 => (x"87",x"d0",x"02",x"98"),
  1277 => (x"48",x"bf",x"d0",x"ff"),
  1278 => (x"98",x"c0",x"c0",x"c8"),
  1279 => (x"70",x"58",x"a6",x"c4"),
  1280 => (x"87",x"f0",x"05",x"98"),
  1281 => (x"c0",x"48",x"d0",x"ff"),
  1282 => (x"1e",x"c7",x"78",x"e0"),
  1283 => (x"e4",x"c1",x"1e",x"c0"),
  1284 => (x"e5",x"c2",x"1e",x"e0"),
  1285 => (x"c1",x"49",x"bf",x"e4"),
  1286 => (x"49",x"74",x"87",x"e1"),
  1287 => (x"87",x"de",x"f7",x"c0"),
  1288 => (x"e7",x"e3",x"8e",x"e4"),
  1289 => (x"1e",x"73",x"1e",x"87"),
  1290 => (x"fc",x"49",x"4b",x"71"),
  1291 => (x"49",x"73",x"87",x"d1"),
  1292 => (x"e3",x"87",x"cc",x"fc"),
  1293 => (x"73",x"1e",x"87",x"da"),
  1294 => (x"c2",x"4b",x"71",x"1e"),
  1295 => (x"d5",x"02",x"4a",x"a3"),
  1296 => (x"05",x"8a",x"c1",x"87"),
  1297 => (x"e5",x"c2",x"87",x"db"),
  1298 => (x"d4",x"02",x"bf",x"f8"),
  1299 => (x"88",x"c1",x"48",x"87"),
  1300 => (x"58",x"fc",x"e5",x"c2"),
  1301 => (x"e5",x"c2",x"87",x"cb"),
  1302 => (x"c1",x"48",x"bf",x"f8"),
  1303 => (x"fc",x"e5",x"c2",x"80"),
  1304 => (x"c0",x"1e",x"c7",x"58"),
  1305 => (x"e0",x"e4",x"c1",x"1e"),
  1306 => (x"e4",x"e5",x"c2",x"1e"),
  1307 => (x"87",x"cb",x"49",x"bf"),
  1308 => (x"f6",x"c0",x"49",x"73"),
  1309 => (x"8e",x"f4",x"87",x"c8"),
  1310 => (x"0e",x"87",x"d5",x"e2"),
  1311 => (x"5d",x"5c",x"5b",x"5e"),
  1312 => (x"86",x"d8",x"ff",x"0e"),
  1313 => (x"c8",x"59",x"a6",x"dc"),
  1314 => (x"78",x"c0",x"48",x"a6"),
  1315 => (x"78",x"c0",x"80",x"c4"),
  1316 => (x"c2",x"80",x"c4",x"4d"),
  1317 => (x"78",x"bf",x"f8",x"e5"),
  1318 => (x"c3",x"48",x"d4",x"ff"),
  1319 => (x"d0",x"ff",x"78",x"ff"),
  1320 => (x"c0",x"c8",x"48",x"bf"),
  1321 => (x"a6",x"c4",x"98",x"c0"),
  1322 => (x"02",x"98",x"70",x"58"),
  1323 => (x"d0",x"ff",x"87",x"d0"),
  1324 => (x"c0",x"c8",x"48",x"bf"),
  1325 => (x"a6",x"c4",x"98",x"c0"),
  1326 => (x"05",x"98",x"70",x"58"),
  1327 => (x"d0",x"ff",x"87",x"f0"),
  1328 => (x"78",x"e1",x"c0",x"48"),
  1329 => (x"d4",x"48",x"d4",x"ff"),
  1330 => (x"f6",x"de",x"ff",x"78"),
  1331 => (x"48",x"d4",x"ff",x"87"),
  1332 => (x"d4",x"78",x"ff",x"c3"),
  1333 => (x"d4",x"ff",x"48",x"a6"),
  1334 => (x"66",x"d4",x"78",x"bf"),
  1335 => (x"a8",x"fb",x"c0",x"48"),
  1336 => (x"87",x"d3",x"c1",x"02"),
  1337 => (x"4a",x"66",x"f8",x"c0"),
  1338 => (x"7e",x"6a",x"82",x"c4"),
  1339 => (x"c2",x"c1",x"1e",x"72"),
  1340 => (x"66",x"c4",x"48",x"f9"),
  1341 => (x"4a",x"a1",x"c8",x"49"),
  1342 => (x"aa",x"71",x"41",x"20"),
  1343 => (x"10",x"87",x"f9",x"05"),
  1344 => (x"c0",x"4a",x"26",x"51"),
  1345 => (x"c8",x"49",x"66",x"f8"),
  1346 => (x"d0",x"cc",x"c1",x"81"),
  1347 => (x"c7",x"49",x"6a",x"79"),
  1348 => (x"51",x"66",x"d4",x"81"),
  1349 => (x"1e",x"d8",x"1e",x"c1"),
  1350 => (x"81",x"c8",x"49",x"6a"),
  1351 => (x"87",x"fa",x"dd",x"ff"),
  1352 => (x"66",x"d0",x"86",x"c8"),
  1353 => (x"a8",x"b7",x"c0",x"48"),
  1354 => (x"c1",x"87",x"c4",x"01"),
  1355 => (x"d0",x"87",x"c8",x"4d"),
  1356 => (x"88",x"c1",x"48",x"66"),
  1357 => (x"d4",x"58",x"a6",x"d4"),
  1358 => (x"f4",x"ca",x"02",x"66"),
  1359 => (x"66",x"c0",x"c1",x"87"),
  1360 => (x"ca",x"03",x"ad",x"b7"),
  1361 => (x"d4",x"ff",x"87",x"eb"),
  1362 => (x"78",x"ff",x"c3",x"48"),
  1363 => (x"ff",x"48",x"a6",x"d4"),
  1364 => (x"d4",x"78",x"bf",x"d4"),
  1365 => (x"c6",x"c1",x"48",x"66"),
  1366 => (x"58",x"a6",x"c4",x"88"),
  1367 => (x"c0",x"02",x"98",x"70"),
  1368 => (x"c9",x"48",x"87",x"e6"),
  1369 => (x"58",x"a6",x"c4",x"88"),
  1370 => (x"c4",x"02",x"98",x"70"),
  1371 => (x"c1",x"48",x"87",x"d5"),
  1372 => (x"58",x"a6",x"c4",x"88"),
  1373 => (x"c1",x"02",x"98",x"70"),
  1374 => (x"c4",x"48",x"87",x"e3"),
  1375 => (x"70",x"58",x"a6",x"88"),
  1376 => (x"fe",x"c3",x"02",x"98"),
  1377 => (x"87",x"d3",x"c9",x"87"),
  1378 => (x"c1",x"05",x"66",x"d8"),
  1379 => (x"d4",x"ff",x"87",x"c5"),
  1380 => (x"78",x"ff",x"c3",x"48"),
  1381 => (x"1e",x"ca",x"1e",x"c0"),
  1382 => (x"93",x"cc",x"4b",x"75"),
  1383 => (x"83",x"66",x"c0",x"c1"),
  1384 => (x"6c",x"4c",x"a3",x"c4"),
  1385 => (x"f1",x"db",x"ff",x"49"),
  1386 => (x"de",x"1e",x"c1",x"87"),
  1387 => (x"ff",x"49",x"6c",x"1e"),
  1388 => (x"d0",x"87",x"e7",x"db"),
  1389 => (x"49",x"a3",x"c8",x"86"),
  1390 => (x"79",x"d0",x"cc",x"c1"),
  1391 => (x"ad",x"b7",x"66",x"d0"),
  1392 => (x"c1",x"87",x"c5",x"04"),
  1393 => (x"87",x"da",x"c8",x"85"),
  1394 => (x"c1",x"48",x"66",x"d0"),
  1395 => (x"58",x"a6",x"d4",x"88"),
  1396 => (x"ff",x"87",x"cf",x"c8"),
  1397 => (x"d8",x"87",x"ec",x"da"),
  1398 => (x"c5",x"c8",x"58",x"a6"),
  1399 => (x"f3",x"dc",x"ff",x"87"),
  1400 => (x"58",x"a6",x"cc",x"87"),
  1401 => (x"a8",x"b7",x"66",x"cc"),
  1402 => (x"cc",x"87",x"c6",x"06"),
  1403 => (x"66",x"c8",x"48",x"a6"),
  1404 => (x"df",x"dc",x"ff",x"78"),
  1405 => (x"a8",x"ec",x"c0",x"87"),
  1406 => (x"87",x"c7",x"c2",x"05"),
  1407 => (x"c1",x"05",x"66",x"d8"),
  1408 => (x"49",x"75",x"87",x"f7"),
  1409 => (x"f8",x"c0",x"91",x"cc"),
  1410 => (x"a1",x"c4",x"81",x"66"),
  1411 => (x"c1",x"4c",x"6a",x"4a"),
  1412 => (x"66",x"c8",x"4a",x"a1"),
  1413 => (x"79",x"97",x"c2",x"52"),
  1414 => (x"cc",x"c1",x"81",x"c8"),
  1415 => (x"d4",x"ff",x"79",x"de"),
  1416 => (x"78",x"ff",x"c3",x"48"),
  1417 => (x"ff",x"48",x"a6",x"d4"),
  1418 => (x"d4",x"78",x"bf",x"d4"),
  1419 => (x"e8",x"c0",x"02",x"66"),
  1420 => (x"fb",x"c0",x"48",x"87"),
  1421 => (x"e0",x"c0",x"02",x"a8"),
  1422 => (x"97",x"66",x"d4",x"87"),
  1423 => (x"ff",x"84",x"c1",x"7c"),
  1424 => (x"ff",x"c3",x"48",x"d4"),
  1425 => (x"48",x"a6",x"d4",x"78"),
  1426 => (x"78",x"bf",x"d4",x"ff"),
  1427 => (x"c8",x"02",x"66",x"d4"),
  1428 => (x"fb",x"c0",x"48",x"87"),
  1429 => (x"e0",x"ff",x"05",x"a8"),
  1430 => (x"54",x"e0",x"c0",x"87"),
  1431 => (x"c0",x"54",x"c1",x"c2"),
  1432 => (x"66",x"d0",x"7c",x"97"),
  1433 => (x"c5",x"04",x"ad",x"b7"),
  1434 => (x"c5",x"85",x"c1",x"87"),
  1435 => (x"66",x"d0",x"87",x"f4"),
  1436 => (x"d4",x"88",x"c1",x"48"),
  1437 => (x"e9",x"c5",x"58",x"a6"),
  1438 => (x"c6",x"d8",x"ff",x"87"),
  1439 => (x"58",x"a6",x"d8",x"87"),
  1440 => (x"c8",x"87",x"df",x"c5"),
  1441 => (x"66",x"d8",x"48",x"66"),
  1442 => (x"c4",x"c5",x"05",x"a8"),
  1443 => (x"48",x"a6",x"dc",x"87"),
  1444 => (x"d9",x"ff",x"78",x"c0"),
  1445 => (x"a6",x"d8",x"87",x"fe"),
  1446 => (x"f7",x"d9",x"ff",x"58"),
  1447 => (x"a6",x"e4",x"c0",x"87"),
  1448 => (x"a8",x"ec",x"c0",x"58"),
  1449 => (x"87",x"ca",x"c0",x"05"),
  1450 => (x"48",x"a6",x"e0",x"c0"),
  1451 => (x"c0",x"78",x"66",x"d4"),
  1452 => (x"d4",x"ff",x"87",x"c6"),
  1453 => (x"78",x"ff",x"c3",x"48"),
  1454 => (x"91",x"cc",x"49",x"75"),
  1455 => (x"48",x"66",x"f8",x"c0"),
  1456 => (x"a6",x"c4",x"80",x"71"),
  1457 => (x"c3",x"49",x"6e",x"58"),
  1458 => (x"51",x"66",x"d4",x"81"),
  1459 => (x"49",x"66",x"e0",x"c0"),
  1460 => (x"66",x"d4",x"81",x"c1"),
  1461 => (x"71",x"48",x"c1",x"89"),
  1462 => (x"c1",x"49",x"70",x"30"),
  1463 => (x"c1",x"4a",x"6e",x"89"),
  1464 => (x"97",x"09",x"72",x"82"),
  1465 => (x"48",x"6e",x"09",x"79"),
  1466 => (x"e5",x"c2",x"50",x"c2"),
  1467 => (x"d4",x"49",x"bf",x"e0"),
  1468 => (x"97",x"29",x"b7",x"66"),
  1469 => (x"71",x"48",x"4a",x"6a"),
  1470 => (x"a6",x"e8",x"c0",x"98"),
  1471 => (x"c4",x"48",x"6e",x"58"),
  1472 => (x"58",x"a6",x"c8",x"80"),
  1473 => (x"4c",x"bf",x"66",x"c4"),
  1474 => (x"c8",x"48",x"66",x"d8"),
  1475 => (x"c0",x"02",x"a8",x"66"),
  1476 => (x"e0",x"c0",x"87",x"c9"),
  1477 => (x"78",x"c0",x"48",x"a6"),
  1478 => (x"c0",x"87",x"c6",x"c0"),
  1479 => (x"c1",x"48",x"a6",x"e0"),
  1480 => (x"66",x"e0",x"c0",x"78"),
  1481 => (x"1e",x"e0",x"c0",x"1e"),
  1482 => (x"d5",x"ff",x"49",x"74"),
  1483 => (x"86",x"c8",x"87",x"ec"),
  1484 => (x"c0",x"58",x"a6",x"d8"),
  1485 => (x"c1",x"06",x"a8",x"b7"),
  1486 => (x"66",x"d4",x"87",x"da"),
  1487 => (x"bf",x"66",x"c4",x"84"),
  1488 => (x"81",x"e0",x"c0",x"49"),
  1489 => (x"c1",x"4b",x"89",x"74"),
  1490 => (x"71",x"4a",x"c2",x"c3"),
  1491 => (x"87",x"e0",x"e5",x"fe"),
  1492 => (x"66",x"dc",x"84",x"c2"),
  1493 => (x"c0",x"80",x"c1",x"48"),
  1494 => (x"c0",x"58",x"a6",x"e0"),
  1495 => (x"c1",x"49",x"66",x"e4"),
  1496 => (x"02",x"a9",x"70",x"81"),
  1497 => (x"c0",x"87",x"c9",x"c0"),
  1498 => (x"c0",x"48",x"a6",x"e0"),
  1499 => (x"87",x"c6",x"c0",x"78"),
  1500 => (x"48",x"a6",x"e0",x"c0"),
  1501 => (x"e0",x"c0",x"78",x"c1"),
  1502 => (x"66",x"c8",x"1e",x"66"),
  1503 => (x"e0",x"c0",x"49",x"bf"),
  1504 => (x"71",x"89",x"74",x"81"),
  1505 => (x"ff",x"49",x"74",x"1e"),
  1506 => (x"c8",x"87",x"cf",x"d4"),
  1507 => (x"a8",x"b7",x"c0",x"86"),
  1508 => (x"87",x"fe",x"fe",x"01"),
  1509 => (x"c0",x"02",x"66",x"dc"),
  1510 => (x"49",x"6e",x"87",x"d2"),
  1511 => (x"66",x"dc",x"81",x"c2"),
  1512 => (x"c8",x"49",x"6e",x"51"),
  1513 => (x"ff",x"cc",x"c1",x"81"),
  1514 => (x"87",x"cd",x"c0",x"79"),
  1515 => (x"81",x"c2",x"49",x"6e"),
  1516 => (x"c8",x"49",x"6e",x"51"),
  1517 => (x"e5",x"d0",x"c1",x"81"),
  1518 => (x"b7",x"66",x"d0",x"79"),
  1519 => (x"c5",x"c0",x"04",x"ad"),
  1520 => (x"c0",x"85",x"c1",x"87"),
  1521 => (x"66",x"d0",x"87",x"dc"),
  1522 => (x"d4",x"88",x"c1",x"48"),
  1523 => (x"d1",x"c0",x"58",x"a6"),
  1524 => (x"ee",x"d2",x"ff",x"87"),
  1525 => (x"58",x"a6",x"d8",x"87"),
  1526 => (x"ff",x"87",x"c7",x"c0"),
  1527 => (x"d8",x"87",x"e4",x"d2"),
  1528 => (x"66",x"d4",x"58",x"a6"),
  1529 => (x"87",x"c9",x"c0",x"02"),
  1530 => (x"b7",x"66",x"c0",x"c1"),
  1531 => (x"d5",x"f5",x"04",x"ad"),
  1532 => (x"ad",x"b7",x"c7",x"87"),
  1533 => (x"87",x"dc",x"c0",x"03"),
  1534 => (x"91",x"cc",x"49",x"75"),
  1535 => (x"81",x"66",x"f8",x"c0"),
  1536 => (x"6a",x"4a",x"a1",x"c4"),
  1537 => (x"c8",x"52",x"c0",x"4a"),
  1538 => (x"c1",x"79",x"c0",x"81"),
  1539 => (x"ad",x"b7",x"c7",x"85"),
  1540 => (x"87",x"e4",x"ff",x"04"),
  1541 => (x"c0",x"02",x"66",x"d8"),
  1542 => (x"f8",x"c0",x"87",x"eb"),
  1543 => (x"d4",x"c1",x"49",x"66"),
  1544 => (x"66",x"f8",x"c0",x"81"),
  1545 => (x"82",x"d5",x"c1",x"4a"),
  1546 => (x"51",x"c2",x"52",x"c0"),
  1547 => (x"49",x"66",x"f8",x"c0"),
  1548 => (x"c1",x"81",x"dc",x"c1"),
  1549 => (x"c0",x"79",x"de",x"cc"),
  1550 => (x"c1",x"49",x"66",x"f8"),
  1551 => (x"c3",x"c1",x"81",x"d8"),
  1552 => (x"d6",x"c0",x"79",x"c5"),
  1553 => (x"66",x"f8",x"c0",x"87"),
  1554 => (x"81",x"d8",x"c1",x"49"),
  1555 => (x"79",x"cc",x"c3",x"c1"),
  1556 => (x"49",x"66",x"f8",x"c0"),
  1557 => (x"c2",x"81",x"dc",x"c1"),
  1558 => (x"c1",x"79",x"f5",x"ca"),
  1559 => (x"c0",x"4a",x"f6",x"d0"),
  1560 => (x"c1",x"49",x"66",x"f8"),
  1561 => (x"79",x"72",x"81",x"e8"),
  1562 => (x"48",x"bf",x"d0",x"ff"),
  1563 => (x"98",x"c0",x"c0",x"c8"),
  1564 => (x"70",x"58",x"a6",x"c4"),
  1565 => (x"d1",x"c0",x"02",x"98"),
  1566 => (x"bf",x"d0",x"ff",x"87"),
  1567 => (x"c0",x"c0",x"c8",x"48"),
  1568 => (x"58",x"a6",x"c4",x"98"),
  1569 => (x"ff",x"05",x"98",x"70"),
  1570 => (x"d0",x"ff",x"87",x"ef"),
  1571 => (x"78",x"e0",x"c0",x"48"),
  1572 => (x"ff",x"48",x"66",x"cc"),
  1573 => (x"d1",x"ff",x"8e",x"d8"),
  1574 => (x"c7",x"1e",x"87",x"f2"),
  1575 => (x"c1",x"1e",x"c0",x"1e"),
  1576 => (x"c2",x"1e",x"e0",x"e4"),
  1577 => (x"49",x"bf",x"e4",x"e5"),
  1578 => (x"c1",x"87",x"d0",x"ef"),
  1579 => (x"c0",x"49",x"e0",x"e4"),
  1580 => (x"f4",x"87",x"e2",x"e7"),
  1581 => (x"1e",x"4f",x"26",x"8e"),
  1582 => (x"c2",x"87",x"c6",x"ca"),
  1583 => (x"c0",x"48",x"c0",x"e6"),
  1584 => (x"48",x"d4",x"ff",x"50"),
  1585 => (x"c1",x"78",x"ff",x"c3"),
  1586 => (x"fe",x"49",x"d3",x"c3"),
  1587 => (x"fe",x"87",x"fd",x"de"),
  1588 => (x"70",x"87",x"c8",x"e8"),
  1589 => (x"87",x"cd",x"02",x"98"),
  1590 => (x"87",x"c5",x"f4",x"fe"),
  1591 => (x"c4",x"02",x"98",x"70"),
  1592 => (x"c2",x"4a",x"c1",x"87"),
  1593 => (x"72",x"4a",x"c0",x"87"),
  1594 => (x"87",x"c8",x"02",x"9a"),
  1595 => (x"49",x"dd",x"c3",x"c1"),
  1596 => (x"87",x"d8",x"de",x"fe"),
  1597 => (x"bf",x"d0",x"d7",x"c2"),
  1598 => (x"e3",x"d5",x"ff",x"49"),
  1599 => (x"f8",x"e5",x"c2",x"87"),
  1600 => (x"c2",x"78",x"c0",x"48"),
  1601 => (x"c0",x"48",x"e4",x"e5"),
  1602 => (x"cd",x"fe",x"49",x"78"),
  1603 => (x"87",x"dd",x"c3",x"87"),
  1604 => (x"c0",x"87",x"c2",x"c9"),
  1605 => (x"ff",x"87",x"ed",x"e6"),
  1606 => (x"4f",x"26",x"87",x"f6"),
  1607 => (x"00",x"00",x"10",x"e0"),
  1608 => (x"00",x"00",x"00",x"02"),
  1609 => (x"00",x"00",x"29",x"90"),
  1610 => (x"00",x"00",x"10",x"42"),
  1611 => (x"00",x"00",x"00",x"02"),
  1612 => (x"00",x"00",x"29",x"ae"),
  1613 => (x"00",x"00",x"10",x"42"),
  1614 => (x"00",x"00",x"00",x"02"),
  1615 => (x"00",x"00",x"29",x"cc"),
  1616 => (x"00",x"00",x"10",x"42"),
  1617 => (x"00",x"00",x"00",x"02"),
  1618 => (x"00",x"00",x"29",x"ea"),
  1619 => (x"00",x"00",x"10",x"42"),
  1620 => (x"00",x"00",x"00",x"02"),
  1621 => (x"00",x"00",x"2a",x"08"),
  1622 => (x"00",x"00",x"10",x"42"),
  1623 => (x"00",x"00",x"00",x"02"),
  1624 => (x"00",x"00",x"2a",x"26"),
  1625 => (x"00",x"00",x"10",x"42"),
  1626 => (x"00",x"00",x"00",x"02"),
  1627 => (x"00",x"00",x"2a",x"44"),
  1628 => (x"00",x"00",x"10",x"42"),
  1629 => (x"00",x"00",x"00",x"02"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"00",x"00",x"13",x"1e"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"11",x"12"),
  1635 => (x"d5",x"c1",x"1e",x"1e"),
  1636 => (x"58",x"a6",x"c4",x"87"),
  1637 => (x"1e",x"4f",x"26",x"26"),
  1638 => (x"f0",x"fe",x"4a",x"71"),
  1639 => (x"cd",x"78",x"c0",x"48"),
  1640 => (x"c1",x"0a",x"7a",x"0a"),
  1641 => (x"fe",x"49",x"ed",x"e6"),
  1642 => (x"26",x"87",x"e1",x"db"),
  1643 => (x"74",x"65",x"53",x"4f"),
  1644 => (x"6e",x"61",x"68",x"20"),
  1645 => (x"72",x"65",x"6c",x"64"),
  1646 => (x"6e",x"49",x"00",x"0a"),
  1647 => (x"74",x"6e",x"69",x"20"),
  1648 => (x"75",x"72",x"72",x"65"),
  1649 => (x"63",x"20",x"74",x"70"),
  1650 => (x"74",x"73",x"6e",x"6f"),
  1651 => (x"74",x"63",x"75",x"72"),
  1652 => (x"00",x"0a",x"72",x"6f"),
  1653 => (x"fa",x"e6",x"c1",x"1e"),
  1654 => (x"ef",x"da",x"fe",x"49"),
  1655 => (x"cc",x"e6",x"c1",x"87"),
  1656 => (x"87",x"f3",x"fe",x"49"),
  1657 => (x"fe",x"1e",x"4f",x"26"),
  1658 => (x"26",x"48",x"bf",x"f0"),
  1659 => (x"f0",x"fe",x"1e",x"4f"),
  1660 => (x"26",x"78",x"c1",x"48"),
  1661 => (x"f0",x"fe",x"1e",x"4f"),
  1662 => (x"26",x"78",x"c0",x"48"),
  1663 => (x"4a",x"71",x"1e",x"4f"),
  1664 => (x"a2",x"c4",x"7a",x"c0"),
  1665 => (x"c8",x"79",x"c0",x"49"),
  1666 => (x"79",x"c0",x"49",x"a2"),
  1667 => (x"c0",x"49",x"a2",x"cc"),
  1668 => (x"0e",x"4f",x"26",x"79"),
  1669 => (x"0e",x"5c",x"5b",x"5e"),
  1670 => (x"4c",x"71",x"86",x"f8"),
  1671 => (x"cc",x"49",x"a4",x"c8"),
  1672 => (x"48",x"6b",x"4b",x"a4"),
  1673 => (x"a6",x"c4",x"80",x"c1"),
  1674 => (x"c8",x"98",x"cf",x"58"),
  1675 => (x"48",x"69",x"58",x"a6"),
  1676 => (x"05",x"a8",x"66",x"c4"),
  1677 => (x"48",x"6b",x"87",x"d4"),
  1678 => (x"a6",x"c4",x"80",x"c1"),
  1679 => (x"c8",x"98",x"cf",x"58"),
  1680 => (x"48",x"69",x"58",x"a6"),
  1681 => (x"02",x"a8",x"66",x"c4"),
  1682 => (x"e8",x"fe",x"87",x"ec"),
  1683 => (x"a4",x"d0",x"c1",x"87"),
  1684 => (x"c4",x"48",x"6b",x"49"),
  1685 => (x"58",x"a6",x"c4",x"90"),
  1686 => (x"66",x"d4",x"81",x"70"),
  1687 => (x"c1",x"48",x"6b",x"79"),
  1688 => (x"58",x"a6",x"c8",x"80"),
  1689 => (x"7b",x"70",x"98",x"cf"),
  1690 => (x"fd",x"87",x"d2",x"c1"),
  1691 => (x"8e",x"f8",x"87",x"ff"),
  1692 => (x"4d",x"26",x"87",x"c2"),
  1693 => (x"4b",x"26",x"4c",x"26"),
  1694 => (x"5e",x"0e",x"4f",x"26"),
  1695 => (x"0e",x"5d",x"5c",x"5b"),
  1696 => (x"4d",x"71",x"86",x"f8"),
  1697 => (x"6d",x"4c",x"a5",x"c4"),
  1698 => (x"05",x"a8",x"6c",x"48"),
  1699 => (x"48",x"ff",x"87",x"c5"),
  1700 => (x"fd",x"87",x"e5",x"c0"),
  1701 => (x"a5",x"d0",x"87",x"df"),
  1702 => (x"c4",x"48",x"6c",x"4b"),
  1703 => (x"58",x"a6",x"c4",x"90"),
  1704 => (x"4b",x"6b",x"83",x"70"),
  1705 => (x"6c",x"9b",x"ff",x"c3"),
  1706 => (x"c8",x"80",x"c1",x"48"),
  1707 => (x"98",x"cf",x"58",x"a6"),
  1708 => (x"f8",x"fc",x"7c",x"70"),
  1709 => (x"48",x"49",x"73",x"87"),
  1710 => (x"f5",x"fe",x"8e",x"f8"),
  1711 => (x"1e",x"73",x"1e",x"87"),
  1712 => (x"f0",x"fc",x"86",x"f8"),
  1713 => (x"4b",x"bf",x"e0",x"87"),
  1714 => (x"c0",x"e0",x"c0",x"49"),
  1715 => (x"e7",x"c0",x"02",x"99"),
  1716 => (x"c3",x"4a",x"73",x"87"),
  1717 => (x"e9",x"c2",x"9a",x"ff"),
  1718 => (x"c4",x"48",x"bf",x"e2"),
  1719 => (x"58",x"a6",x"c4",x"90"),
  1720 => (x"49",x"f2",x"e9",x"c2"),
  1721 => (x"79",x"72",x"81",x"70"),
  1722 => (x"bf",x"e2",x"e9",x"c2"),
  1723 => (x"c8",x"80",x"c1",x"48"),
  1724 => (x"98",x"cf",x"58",x"a6"),
  1725 => (x"58",x"e6",x"e9",x"c2"),
  1726 => (x"c0",x"d0",x"49",x"73"),
  1727 => (x"f2",x"c0",x"02",x"99"),
  1728 => (x"ea",x"e9",x"c2",x"87"),
  1729 => (x"e9",x"c2",x"48",x"bf"),
  1730 => (x"02",x"a8",x"bf",x"ee"),
  1731 => (x"c2",x"87",x"e4",x"c0"),
  1732 => (x"48",x"bf",x"ea",x"e9"),
  1733 => (x"a6",x"c4",x"90",x"c4"),
  1734 => (x"f2",x"ea",x"c2",x"58"),
  1735 => (x"e0",x"81",x"70",x"49"),
  1736 => (x"c2",x"78",x"69",x"48"),
  1737 => (x"48",x"bf",x"ea",x"e9"),
  1738 => (x"a6",x"c8",x"80",x"c1"),
  1739 => (x"c2",x"98",x"cf",x"58"),
  1740 => (x"fa",x"58",x"ee",x"e9"),
  1741 => (x"a6",x"c4",x"87",x"f0"),
  1742 => (x"87",x"f1",x"fa",x"58"),
  1743 => (x"f5",x"fc",x"8e",x"f8"),
  1744 => (x"e9",x"c2",x"1e",x"87"),
  1745 => (x"f4",x"fa",x"49",x"e2"),
  1746 => (x"fd",x"ea",x"c1",x"87"),
  1747 => (x"87",x"c7",x"f9",x"49"),
  1748 => (x"26",x"87",x"f5",x"c3"),
  1749 => (x"1e",x"73",x"1e",x"4f"),
  1750 => (x"49",x"e2",x"e9",x"c2"),
  1751 => (x"70",x"87",x"db",x"fc"),
  1752 => (x"aa",x"b7",x"c0",x"4a"),
  1753 => (x"87",x"cc",x"c2",x"04"),
  1754 => (x"05",x"aa",x"f0",x"c3"),
  1755 => (x"f0",x"c1",x"87",x"c9"),
  1756 => (x"78",x"c1",x"48",x"c0"),
  1757 => (x"c3",x"87",x"ed",x"c1"),
  1758 => (x"c9",x"05",x"aa",x"e0"),
  1759 => (x"c4",x"f0",x"c1",x"87"),
  1760 => (x"c1",x"78",x"c1",x"48"),
  1761 => (x"f0",x"c1",x"87",x"de"),
  1762 => (x"c6",x"02",x"bf",x"c4"),
  1763 => (x"a2",x"c0",x"c2",x"87"),
  1764 => (x"72",x"87",x"c2",x"4b"),
  1765 => (x"c0",x"f0",x"c1",x"4b"),
  1766 => (x"e0",x"c0",x"02",x"bf"),
  1767 => (x"c4",x"49",x"73",x"87"),
  1768 => (x"c1",x"91",x"29",x"b7"),
  1769 => (x"73",x"81",x"c8",x"f0"),
  1770 => (x"c2",x"9a",x"cf",x"4a"),
  1771 => (x"72",x"48",x"c1",x"92"),
  1772 => (x"ff",x"4a",x"70",x"30"),
  1773 => (x"69",x"48",x"72",x"ba"),
  1774 => (x"db",x"79",x"70",x"98"),
  1775 => (x"c4",x"49",x"73",x"87"),
  1776 => (x"c1",x"91",x"29",x"b7"),
  1777 => (x"73",x"81",x"c8",x"f0"),
  1778 => (x"c2",x"9a",x"cf",x"4a"),
  1779 => (x"72",x"48",x"c3",x"92"),
  1780 => (x"48",x"4a",x"70",x"30"),
  1781 => (x"79",x"70",x"b0",x"69"),
  1782 => (x"48",x"c4",x"f0",x"c1"),
  1783 => (x"f0",x"c1",x"78",x"c0"),
  1784 => (x"78",x"c0",x"48",x"c0"),
  1785 => (x"49",x"e2",x"e9",x"c2"),
  1786 => (x"70",x"87",x"cf",x"fa"),
  1787 => (x"aa",x"b7",x"c0",x"4a"),
  1788 => (x"87",x"f4",x"fd",x"03"),
  1789 => (x"87",x"c4",x"48",x"c0"),
  1790 => (x"4c",x"26",x"4d",x"26"),
  1791 => (x"4f",x"26",x"4b",x"26"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"00",x"00",x"00",x"00"),
  1807 => (x"00",x"00",x"00",x"00"),
  1808 => (x"00",x"00",x"00",x"00"),
  1809 => (x"00",x"00",x"00",x"00"),
  1810 => (x"72",x"4a",x"c0",x"1e"),
  1811 => (x"c1",x"91",x"c4",x"49"),
  1812 => (x"c0",x"81",x"c8",x"f0"),
  1813 => (x"d0",x"82",x"c1",x"79"),
  1814 => (x"ee",x"04",x"aa",x"b7"),
  1815 => (x"0e",x"4f",x"26",x"87"),
  1816 => (x"5d",x"5c",x"5b",x"5e"),
  1817 => (x"f6",x"4d",x"71",x"0e"),
  1818 => (x"4a",x"75",x"87",x"cb"),
  1819 => (x"92",x"2a",x"b7",x"c4"),
  1820 => (x"82",x"c8",x"f0",x"c1"),
  1821 => (x"9c",x"cf",x"4c",x"75"),
  1822 => (x"49",x"6a",x"94",x"c2"),
  1823 => (x"c3",x"2b",x"74",x"4b"),
  1824 => (x"74",x"48",x"c2",x"9b"),
  1825 => (x"ff",x"4c",x"70",x"30"),
  1826 => (x"71",x"48",x"74",x"bc"),
  1827 => (x"f5",x"7a",x"70",x"98"),
  1828 => (x"48",x"73",x"87",x"db"),
  1829 => (x"1e",x"87",x"e1",x"fd"),
  1830 => (x"bf",x"d0",x"ff",x"1e"),
  1831 => (x"c0",x"c0",x"c8",x"48"),
  1832 => (x"58",x"a6",x"c4",x"98"),
  1833 => (x"d0",x"02",x"98",x"70"),
  1834 => (x"bf",x"d0",x"ff",x"87"),
  1835 => (x"c0",x"c0",x"c8",x"48"),
  1836 => (x"58",x"a6",x"c4",x"98"),
  1837 => (x"f0",x"05",x"98",x"70"),
  1838 => (x"48",x"d0",x"ff",x"87"),
  1839 => (x"71",x"78",x"e1",x"c4"),
  1840 => (x"08",x"d4",x"ff",x"48"),
  1841 => (x"48",x"66",x"c8",x"78"),
  1842 => (x"78",x"08",x"d4",x"ff"),
  1843 => (x"1e",x"4f",x"26",x"26"),
  1844 => (x"c8",x"4a",x"71",x"1e"),
  1845 => (x"72",x"1e",x"49",x"66"),
  1846 => (x"87",x"fb",x"fe",x"49"),
  1847 => (x"d0",x"ff",x"86",x"c4"),
  1848 => (x"c0",x"c8",x"48",x"bf"),
  1849 => (x"a6",x"c4",x"98",x"c0"),
  1850 => (x"02",x"98",x"70",x"58"),
  1851 => (x"d0",x"ff",x"87",x"d0"),
  1852 => (x"c0",x"c8",x"48",x"bf"),
  1853 => (x"a6",x"c4",x"98",x"c0"),
  1854 => (x"05",x"98",x"70",x"58"),
  1855 => (x"d0",x"ff",x"87",x"f0"),
  1856 => (x"78",x"e0",x"c0",x"48"),
  1857 => (x"1e",x"4f",x"26",x"26"),
  1858 => (x"4b",x"71",x"1e",x"73"),
  1859 => (x"73",x"1e",x"66",x"c8"),
  1860 => (x"a2",x"e0",x"c1",x"4a"),
  1861 => (x"87",x"f7",x"fe",x"49"),
  1862 => (x"26",x"87",x"c4",x"26"),
  1863 => (x"26",x"4c",x"26",x"4d"),
  1864 => (x"1e",x"4f",x"26",x"4b"),
  1865 => (x"bf",x"d0",x"ff",x"1e"),
  1866 => (x"c0",x"c0",x"c8",x"48"),
  1867 => (x"58",x"a6",x"c4",x"98"),
  1868 => (x"d0",x"02",x"98",x"70"),
  1869 => (x"bf",x"d0",x"ff",x"87"),
  1870 => (x"c0",x"c0",x"c8",x"48"),
  1871 => (x"58",x"a6",x"c4",x"98"),
  1872 => (x"f0",x"05",x"98",x"70"),
  1873 => (x"48",x"d0",x"ff",x"87"),
  1874 => (x"71",x"78",x"c9",x"c4"),
  1875 => (x"08",x"d4",x"ff",x"48"),
  1876 => (x"4f",x"26",x"26",x"78"),
  1877 => (x"4a",x"71",x"1e",x"1e"),
  1878 => (x"87",x"c7",x"ff",x"49"),
  1879 => (x"48",x"bf",x"d0",x"ff"),
  1880 => (x"98",x"c0",x"c0",x"c8"),
  1881 => (x"70",x"58",x"a6",x"c4"),
  1882 => (x"87",x"d0",x"02",x"98"),
  1883 => (x"48",x"bf",x"d0",x"ff"),
  1884 => (x"98",x"c0",x"c0",x"c8"),
  1885 => (x"70",x"58",x"a6",x"c4"),
  1886 => (x"87",x"f0",x"05",x"98"),
  1887 => (x"c8",x"48",x"d0",x"ff"),
  1888 => (x"4f",x"26",x"26",x"78"),
  1889 => (x"1e",x"1e",x"73",x"1e"),
  1890 => (x"eb",x"c2",x"4b",x"71"),
  1891 => (x"c3",x"02",x"bf",x"fe"),
  1892 => (x"87",x"cc",x"c3",x"87"),
  1893 => (x"48",x"bf",x"d0",x"ff"),
  1894 => (x"98",x"c0",x"c0",x"c8"),
  1895 => (x"70",x"58",x"a6",x"c4"),
  1896 => (x"87",x"d0",x"02",x"98"),
  1897 => (x"48",x"bf",x"d0",x"ff"),
  1898 => (x"98",x"c0",x"c0",x"c8"),
  1899 => (x"70",x"58",x"a6",x"c4"),
  1900 => (x"87",x"f0",x"05",x"98"),
  1901 => (x"c4",x"48",x"d0",x"ff"),
  1902 => (x"48",x"73",x"78",x"c9"),
  1903 => (x"ff",x"b0",x"e0",x"c0"),
  1904 => (x"c2",x"78",x"08",x"d4"),
  1905 => (x"c0",x"48",x"f2",x"eb"),
  1906 => (x"02",x"66",x"cc",x"78"),
  1907 => (x"ff",x"c3",x"87",x"c5"),
  1908 => (x"c0",x"87",x"c2",x"49"),
  1909 => (x"fa",x"eb",x"c2",x"49"),
  1910 => (x"02",x"66",x"d0",x"59"),
  1911 => (x"d5",x"c5",x"87",x"c6"),
  1912 => (x"87",x"c4",x"4a",x"d5"),
  1913 => (x"4a",x"ff",x"ff",x"cf"),
  1914 => (x"5a",x"fe",x"eb",x"c2"),
  1915 => (x"48",x"fe",x"eb",x"c2"),
  1916 => (x"c4",x"26",x"78",x"c1"),
  1917 => (x"26",x"4d",x"26",x"87"),
  1918 => (x"26",x"4b",x"26",x"4c"),
  1919 => (x"5b",x"5e",x"0e",x"4f"),
  1920 => (x"71",x"0e",x"5d",x"5c"),
  1921 => (x"fa",x"eb",x"c2",x"4a"),
  1922 => (x"9a",x"72",x"4c",x"bf"),
  1923 => (x"49",x"87",x"cb",x"02"),
  1924 => (x"f6",x"c1",x"91",x"c8"),
  1925 => (x"83",x"71",x"4b",x"fe"),
  1926 => (x"fa",x"c1",x"87",x"c4"),
  1927 => (x"4d",x"c0",x"4b",x"fe"),
  1928 => (x"99",x"74",x"49",x"13"),
  1929 => (x"bf",x"f6",x"eb",x"c2"),
  1930 => (x"ff",x"b8",x"71",x"48"),
  1931 => (x"c1",x"78",x"08",x"d4"),
  1932 => (x"c8",x"85",x"2c",x"b7"),
  1933 => (x"e7",x"04",x"ad",x"b7"),
  1934 => (x"f2",x"eb",x"c2",x"87"),
  1935 => (x"80",x"c8",x"48",x"bf"),
  1936 => (x"58",x"f6",x"eb",x"c2"),
  1937 => (x"1e",x"87",x"ee",x"fe"),
  1938 => (x"4b",x"71",x"1e",x"73"),
  1939 => (x"02",x"9a",x"4a",x"13"),
  1940 => (x"49",x"72",x"87",x"cb"),
  1941 => (x"13",x"87",x"e6",x"fe"),
  1942 => (x"f5",x"05",x"9a",x"4a"),
  1943 => (x"87",x"d9",x"fe",x"87"),
  1944 => (x"eb",x"c2",x"1e",x"1e"),
  1945 => (x"c2",x"49",x"bf",x"f2"),
  1946 => (x"c1",x"48",x"f2",x"eb"),
  1947 => (x"c0",x"c4",x"78",x"a1"),
  1948 => (x"db",x"03",x"a9",x"b7"),
  1949 => (x"48",x"d4",x"ff",x"87"),
  1950 => (x"bf",x"f6",x"eb",x"c2"),
  1951 => (x"f2",x"eb",x"c2",x"78"),
  1952 => (x"eb",x"c2",x"49",x"bf"),
  1953 => (x"a1",x"c1",x"48",x"f2"),
  1954 => (x"b7",x"c0",x"c4",x"78"),
  1955 => (x"87",x"e5",x"04",x"a9"),
  1956 => (x"48",x"bf",x"d0",x"ff"),
  1957 => (x"98",x"c0",x"c0",x"c8"),
  1958 => (x"70",x"58",x"a6",x"c4"),
  1959 => (x"87",x"d0",x"02",x"98"),
  1960 => (x"48",x"bf",x"d0",x"ff"),
  1961 => (x"98",x"c0",x"c0",x"c8"),
  1962 => (x"70",x"58",x"a6",x"c4"),
  1963 => (x"87",x"f0",x"05",x"98"),
  1964 => (x"c8",x"48",x"d0",x"ff"),
  1965 => (x"fe",x"eb",x"c2",x"78"),
  1966 => (x"26",x"78",x"c0",x"48"),
  1967 => (x"00",x"00",x"4f",x"26"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"00",x"00",x"00"),
  1970 => (x"00",x"5f",x"5f",x"00"),
  1971 => (x"03",x"00",x"00",x"00"),
  1972 => (x"03",x"03",x"00",x"03"),
  1973 => (x"7f",x"14",x"00",x"00"),
  1974 => (x"7f",x"7f",x"14",x"7f"),
  1975 => (x"24",x"00",x"00",x"14"),
  1976 => (x"3a",x"6b",x"6b",x"2e"),
  1977 => (x"6a",x"4c",x"00",x"12"),
  1978 => (x"56",x"6c",x"18",x"36"),
  1979 => (x"7e",x"30",x"00",x"32"),
  1980 => (x"3a",x"77",x"59",x"4f"),
  1981 => (x"00",x"00",x"40",x"68"),
  1982 => (x"00",x"03",x"07",x"04"),
  1983 => (x"00",x"00",x"00",x"00"),
  1984 => (x"41",x"63",x"3e",x"1c"),
  1985 => (x"00",x"00",x"00",x"00"),
  1986 => (x"1c",x"3e",x"63",x"41"),
  1987 => (x"2a",x"08",x"00",x"00"),
  1988 => (x"3e",x"1c",x"1c",x"3e"),
  1989 => (x"08",x"00",x"08",x"2a"),
  1990 => (x"08",x"3e",x"3e",x"08"),
  1991 => (x"00",x"00",x"00",x"08"),
  1992 => (x"00",x"60",x"e0",x"80"),
  1993 => (x"08",x"00",x"00",x"00"),
  1994 => (x"08",x"08",x"08",x"08"),
  1995 => (x"00",x"00",x"00",x"08"),
  1996 => (x"00",x"60",x"60",x"00"),
  1997 => (x"60",x"40",x"00",x"00"),
  1998 => (x"06",x"0c",x"18",x"30"),
  1999 => (x"3e",x"00",x"01",x"03"),
  2000 => (x"7f",x"4d",x"59",x"7f"),
  2001 => (x"04",x"00",x"00",x"3e"),
  2002 => (x"00",x"7f",x"7f",x"06"),
  2003 => (x"42",x"00",x"00",x"00"),
  2004 => (x"4f",x"59",x"71",x"63"),
  2005 => (x"22",x"00",x"00",x"46"),
  2006 => (x"7f",x"49",x"49",x"63"),
  2007 => (x"1c",x"18",x"00",x"36"),
  2008 => (x"7f",x"7f",x"13",x"16"),
  2009 => (x"27",x"00",x"00",x"10"),
  2010 => (x"7d",x"45",x"45",x"67"),
  2011 => (x"3c",x"00",x"00",x"39"),
  2012 => (x"79",x"49",x"4b",x"7e"),
  2013 => (x"01",x"00",x"00",x"30"),
  2014 => (x"0f",x"79",x"71",x"01"),
  2015 => (x"36",x"00",x"00",x"07"),
  2016 => (x"7f",x"49",x"49",x"7f"),
  2017 => (x"06",x"00",x"00",x"36"),
  2018 => (x"3f",x"69",x"49",x"4f"),
  2019 => (x"00",x"00",x"00",x"1e"),
  2020 => (x"00",x"66",x"66",x"00"),
  2021 => (x"00",x"00",x"00",x"00"),
  2022 => (x"00",x"66",x"e6",x"80"),
  2023 => (x"08",x"00",x"00",x"00"),
  2024 => (x"22",x"14",x"14",x"08"),
  2025 => (x"14",x"00",x"00",x"22"),
  2026 => (x"14",x"14",x"14",x"14"),
  2027 => (x"22",x"00",x"00",x"14"),
  2028 => (x"08",x"14",x"14",x"22"),
  2029 => (x"02",x"00",x"00",x"08"),
  2030 => (x"0f",x"59",x"51",x"03"),
  2031 => (x"7f",x"3e",x"00",x"06"),
  2032 => (x"1f",x"55",x"5d",x"41"),
  2033 => (x"7e",x"00",x"00",x"1e"),
  2034 => (x"7f",x"09",x"09",x"7f"),
  2035 => (x"7f",x"00",x"00",x"7e"),
  2036 => (x"7f",x"49",x"49",x"7f"),
  2037 => (x"1c",x"00",x"00",x"36"),
  2038 => (x"41",x"41",x"63",x"3e"),
  2039 => (x"7f",x"00",x"00",x"41"),
  2040 => (x"3e",x"63",x"41",x"7f"),
  2041 => (x"7f",x"00",x"00",x"1c"),
  2042 => (x"41",x"49",x"49",x"7f"),
  2043 => (x"7f",x"00",x"00",x"41"),
  2044 => (x"01",x"09",x"09",x"7f"),
  2045 => (x"3e",x"00",x"00",x"01"),
  2046 => (x"7b",x"49",x"41",x"7f"),
  2047 => (x"7f",x"00",x"00",x"7a"),
  2048 => (x"7f",x"08",x"08",x"7f"),
  2049 => (x"00",x"00",x"00",x"7f"),
  2050 => (x"41",x"7f",x"7f",x"41"),
  2051 => (x"20",x"00",x"00",x"00"),
  2052 => (x"7f",x"40",x"40",x"60"),
  2053 => (x"7f",x"7f",x"00",x"3f"),
  2054 => (x"63",x"36",x"1c",x"08"),
  2055 => (x"7f",x"00",x"00",x"41"),
  2056 => (x"40",x"40",x"40",x"7f"),
  2057 => (x"7f",x"7f",x"00",x"40"),
  2058 => (x"7f",x"06",x"0c",x"06"),
  2059 => (x"7f",x"7f",x"00",x"7f"),
  2060 => (x"7f",x"18",x"0c",x"06"),
  2061 => (x"3e",x"00",x"00",x"7f"),
  2062 => (x"7f",x"41",x"41",x"7f"),
  2063 => (x"7f",x"00",x"00",x"3e"),
  2064 => (x"0f",x"09",x"09",x"7f"),
  2065 => (x"7f",x"3e",x"00",x"06"),
  2066 => (x"7e",x"7f",x"61",x"41"),
  2067 => (x"7f",x"00",x"00",x"40"),
  2068 => (x"7f",x"19",x"09",x"7f"),
  2069 => (x"26",x"00",x"00",x"66"),
  2070 => (x"7b",x"59",x"4d",x"6f"),
  2071 => (x"01",x"00",x"00",x"32"),
  2072 => (x"01",x"7f",x"7f",x"01"),
  2073 => (x"3f",x"00",x"00",x"01"),
  2074 => (x"7f",x"40",x"40",x"7f"),
  2075 => (x"0f",x"00",x"00",x"3f"),
  2076 => (x"3f",x"70",x"70",x"3f"),
  2077 => (x"7f",x"7f",x"00",x"0f"),
  2078 => (x"7f",x"30",x"18",x"30"),
  2079 => (x"63",x"41",x"00",x"7f"),
  2080 => (x"36",x"1c",x"1c",x"36"),
  2081 => (x"03",x"01",x"41",x"63"),
  2082 => (x"06",x"7c",x"7c",x"06"),
  2083 => (x"71",x"61",x"01",x"03"),
  2084 => (x"43",x"47",x"4d",x"59"),
  2085 => (x"00",x"00",x"00",x"41"),
  2086 => (x"41",x"41",x"7f",x"7f"),
  2087 => (x"03",x"01",x"00",x"00"),
  2088 => (x"30",x"18",x"0c",x"06"),
  2089 => (x"00",x"00",x"40",x"60"),
  2090 => (x"7f",x"7f",x"41",x"41"),
  2091 => (x"0c",x"08",x"00",x"00"),
  2092 => (x"0c",x"06",x"03",x"06"),
  2093 => (x"80",x"80",x"00",x"08"),
  2094 => (x"80",x"80",x"80",x"80"),
  2095 => (x"00",x"00",x"00",x"80"),
  2096 => (x"04",x"07",x"03",x"00"),
  2097 => (x"20",x"00",x"00",x"00"),
  2098 => (x"7c",x"54",x"54",x"74"),
  2099 => (x"7f",x"00",x"00",x"78"),
  2100 => (x"7c",x"44",x"44",x"7f"),
  2101 => (x"38",x"00",x"00",x"38"),
  2102 => (x"44",x"44",x"44",x"7c"),
  2103 => (x"38",x"00",x"00",x"00"),
  2104 => (x"7f",x"44",x"44",x"7c"),
  2105 => (x"38",x"00",x"00",x"7f"),
  2106 => (x"5c",x"54",x"54",x"7c"),
  2107 => (x"04",x"00",x"00",x"18"),
  2108 => (x"05",x"05",x"7f",x"7e"),
  2109 => (x"18",x"00",x"00",x"00"),
  2110 => (x"fc",x"a4",x"a4",x"bc"),
  2111 => (x"7f",x"00",x"00",x"7c"),
  2112 => (x"7c",x"04",x"04",x"7f"),
  2113 => (x"00",x"00",x"00",x"78"),
  2114 => (x"40",x"7d",x"3d",x"00"),
  2115 => (x"80",x"00",x"00",x"00"),
  2116 => (x"7d",x"fd",x"80",x"80"),
  2117 => (x"7f",x"00",x"00",x"00"),
  2118 => (x"6c",x"38",x"10",x"7f"),
  2119 => (x"00",x"00",x"00",x"44"),
  2120 => (x"40",x"7f",x"3f",x"00"),
  2121 => (x"7c",x"7c",x"00",x"00"),
  2122 => (x"7c",x"0c",x"18",x"0c"),
  2123 => (x"7c",x"00",x"00",x"78"),
  2124 => (x"7c",x"04",x"04",x"7c"),
  2125 => (x"38",x"00",x"00",x"78"),
  2126 => (x"7c",x"44",x"44",x"7c"),
  2127 => (x"fc",x"00",x"00",x"38"),
  2128 => (x"3c",x"24",x"24",x"fc"),
  2129 => (x"18",x"00",x"00",x"18"),
  2130 => (x"fc",x"24",x"24",x"3c"),
  2131 => (x"7c",x"00",x"00",x"fc"),
  2132 => (x"0c",x"04",x"04",x"7c"),
  2133 => (x"48",x"00",x"00",x"08"),
  2134 => (x"74",x"54",x"54",x"5c"),
  2135 => (x"04",x"00",x"00",x"20"),
  2136 => (x"44",x"44",x"7f",x"3f"),
  2137 => (x"3c",x"00",x"00",x"00"),
  2138 => (x"7c",x"40",x"40",x"7c"),
  2139 => (x"1c",x"00",x"00",x"7c"),
  2140 => (x"3c",x"60",x"60",x"3c"),
  2141 => (x"7c",x"3c",x"00",x"1c"),
  2142 => (x"7c",x"60",x"30",x"60"),
  2143 => (x"6c",x"44",x"00",x"3c"),
  2144 => (x"6c",x"38",x"10",x"38"),
  2145 => (x"1c",x"00",x"00",x"44"),
  2146 => (x"3c",x"60",x"e0",x"bc"),
  2147 => (x"44",x"00",x"00",x"1c"),
  2148 => (x"4c",x"5c",x"74",x"64"),
  2149 => (x"08",x"00",x"00",x"44"),
  2150 => (x"41",x"77",x"3e",x"08"),
  2151 => (x"00",x"00",x"00",x"41"),
  2152 => (x"00",x"7f",x"7f",x"00"),
  2153 => (x"41",x"00",x"00",x"00"),
  2154 => (x"08",x"3e",x"77",x"41"),
  2155 => (x"01",x"02",x"00",x"08"),
  2156 => (x"02",x"02",x"03",x"01"),
  2157 => (x"7f",x"7f",x"00",x"01"),
  2158 => (x"7f",x"7f",x"7f",x"7f"),
  2159 => (x"08",x"08",x"00",x"7f"),
  2160 => (x"3e",x"3e",x"1c",x"1c"),
  2161 => (x"7f",x"7f",x"7f",x"7f"),
  2162 => (x"1c",x"1c",x"3e",x"3e"),
  2163 => (x"10",x"00",x"08",x"08"),
  2164 => (x"18",x"7c",x"7c",x"18"),
  2165 => (x"10",x"00",x"00",x"10"),
  2166 => (x"30",x"7c",x"7c",x"30"),
  2167 => (x"30",x"10",x"00",x"10"),
  2168 => (x"1e",x"78",x"60",x"60"),
  2169 => (x"66",x"42",x"00",x"06"),
  2170 => (x"66",x"3c",x"18",x"3c"),
  2171 => (x"38",x"78",x"00",x"42"),
  2172 => (x"6c",x"c6",x"c2",x"6a"),
  2173 => (x"00",x"60",x"00",x"38"),
  2174 => (x"00",x"00",x"60",x"00"),
  2175 => (x"5e",x"0e",x"00",x"60"),
  2176 => (x"0e",x"5d",x"5c",x"5b"),
  2177 => (x"c2",x"4c",x"71",x"1e"),
  2178 => (x"4b",x"bf",x"c6",x"ec"),
  2179 => (x"48",x"ca",x"ec",x"c2"),
  2180 => (x"06",x"27",x"78",x"c0"),
  2181 => (x"bf",x"00",x"00",x"2b"),
  2182 => (x"99",x"49",x"bf",x"97"),
  2183 => (x"87",x"c8",x"c1",x"02"),
  2184 => (x"ec",x"c2",x"1e",x"c0"),
  2185 => (x"74",x"4d",x"bf",x"ca"),
  2186 => (x"87",x"c7",x"02",x"ad"),
  2187 => (x"c0",x"48",x"a6",x"c4"),
  2188 => (x"c4",x"87",x"c5",x"78"),
  2189 => (x"78",x"c1",x"48",x"a6"),
  2190 => (x"75",x"1e",x"66",x"c4"),
  2191 => (x"87",x"c4",x"ed",x"49"),
  2192 => (x"e0",x"c0",x"86",x"c8"),
  2193 => (x"87",x"f5",x"ee",x"49"),
  2194 => (x"6a",x"4a",x"a3",x"c4"),
  2195 => (x"87",x"f7",x"ef",x"49"),
  2196 => (x"c2",x"87",x"cd",x"f0"),
  2197 => (x"48",x"bf",x"ca",x"ec"),
  2198 => (x"ec",x"c2",x"80",x"c1"),
  2199 => (x"83",x"cc",x"58",x"ce"),
  2200 => (x"99",x"49",x"6b",x"97"),
  2201 => (x"87",x"f8",x"fe",x"05"),
  2202 => (x"bf",x"ca",x"ec",x"c2"),
  2203 => (x"ad",x"b7",x"c8",x"4d"),
  2204 => (x"c0",x"87",x"d9",x"03"),
  2205 => (x"ec",x"c2",x"1e",x"1e"),
  2206 => (x"ec",x"49",x"bf",x"ca"),
  2207 => (x"86",x"c8",x"87",x"c6"),
  2208 => (x"c1",x"87",x"dd",x"ef"),
  2209 => (x"ad",x"b7",x"c8",x"85"),
  2210 => (x"87",x"e7",x"ff",x"04"),
  2211 => (x"26",x"4d",x"26",x"26"),
  2212 => (x"26",x"4b",x"26",x"4c"),
  2213 => (x"4a",x"71",x"1e",x"4f"),
  2214 => (x"5a",x"ca",x"ec",x"c2"),
  2215 => (x"bf",x"ce",x"ec",x"c2"),
  2216 => (x"87",x"da",x"fd",x"49"),
  2217 => (x"bf",x"ca",x"ec",x"c2"),
  2218 => (x"c2",x"89",x"c1",x"49"),
  2219 => (x"71",x"59",x"d2",x"ec"),
  2220 => (x"26",x"87",x"cb",x"fd"),
  2221 => (x"c0",x"c1",x"1e",x"4f"),
  2222 => (x"87",x"d8",x"ea",x"49"),
  2223 => (x"48",x"fb",x"d6",x"c2"),
  2224 => (x"4f",x"26",x"78",x"c0"),
  2225 => (x"5c",x"5b",x"5e",x"0e"),
  2226 => (x"86",x"f4",x"0e",x"5d"),
  2227 => (x"c0",x"48",x"a6",x"c8"),
  2228 => (x"7e",x"bf",x"ec",x"78"),
  2229 => (x"ec",x"c2",x"80",x"fc"),
  2230 => (x"c2",x"78",x"bf",x"c6"),
  2231 => (x"4d",x"bf",x"d2",x"ec"),
  2232 => (x"c7",x"4c",x"bf",x"e8"),
  2233 => (x"87",x"f7",x"e5",x"49"),
  2234 => (x"99",x"c2",x"49",x"70"),
  2235 => (x"c2",x"87",x"cf",x"05"),
  2236 => (x"49",x"bf",x"f3",x"d6"),
  2237 => (x"99",x"6e",x"b9",x"ff"),
  2238 => (x"c0",x"02",x"99",x"c1"),
  2239 => (x"49",x"c7",x"87",x"ee"),
  2240 => (x"70",x"87",x"dc",x"e5"),
  2241 => (x"87",x"cd",x"02",x"98"),
  2242 => (x"c7",x"87",x"ca",x"e1"),
  2243 => (x"87",x"cf",x"e5",x"49"),
  2244 => (x"f3",x"05",x"98",x"70"),
  2245 => (x"fb",x"d6",x"c2",x"87"),
  2246 => (x"ba",x"c1",x"4a",x"bf"),
  2247 => (x"5a",x"ff",x"d6",x"c2"),
  2248 => (x"49",x"a2",x"c0",x"c1"),
  2249 => (x"c8",x"87",x"ed",x"e8"),
  2250 => (x"78",x"c1",x"48",x"a6"),
  2251 => (x"48",x"f3",x"d6",x"c2"),
  2252 => (x"d6",x"c2",x"78",x"6e"),
  2253 => (x"c1",x"05",x"bf",x"fb"),
  2254 => (x"a6",x"c4",x"87",x"da"),
  2255 => (x"c0",x"c0",x"c8",x"48"),
  2256 => (x"ff",x"d6",x"c2",x"78"),
  2257 => (x"bf",x"97",x"6e",x"7e"),
  2258 => (x"c1",x"48",x"6e",x"49"),
  2259 => (x"58",x"a6",x"c4",x"80"),
  2260 => (x"87",x"cb",x"e4",x"71"),
  2261 => (x"c3",x"02",x"98",x"70"),
  2262 => (x"b4",x"66",x"c4",x"87"),
  2263 => (x"c1",x"48",x"66",x"c4"),
  2264 => (x"a6",x"c8",x"28",x"b7"),
  2265 => (x"05",x"98",x"70",x"58"),
  2266 => (x"74",x"87",x"da",x"ff"),
  2267 => (x"99",x"ff",x"c3",x"49"),
  2268 => (x"49",x"c0",x"1e",x"71"),
  2269 => (x"74",x"87",x"d0",x"e6"),
  2270 => (x"29",x"b7",x"c8",x"49"),
  2271 => (x"49",x"c1",x"1e",x"71"),
  2272 => (x"c8",x"87",x"c4",x"e6"),
  2273 => (x"49",x"fd",x"c3",x"86"),
  2274 => (x"c3",x"87",x"d4",x"e3"),
  2275 => (x"ce",x"e3",x"49",x"fa"),
  2276 => (x"87",x"ca",x"c8",x"87"),
  2277 => (x"ff",x"c3",x"49",x"74"),
  2278 => (x"2c",x"b7",x"c8",x"99"),
  2279 => (x"9c",x"74",x"b4",x"71"),
  2280 => (x"ff",x"87",x"dd",x"02"),
  2281 => (x"6e",x"7e",x"bf",x"c8"),
  2282 => (x"f7",x"d6",x"c2",x"49"),
  2283 => (x"c0",x"c2",x"89",x"bf"),
  2284 => (x"87",x"c4",x"03",x"a9"),
  2285 => (x"87",x"ce",x"4c",x"c0"),
  2286 => (x"48",x"f7",x"d6",x"c2"),
  2287 => (x"87",x"c6",x"78",x"6e"),
  2288 => (x"48",x"f7",x"d6",x"c2"),
  2289 => (x"49",x"74",x"78",x"c0"),
  2290 => (x"ce",x"05",x"99",x"c8"),
  2291 => (x"49",x"f5",x"c3",x"87"),
  2292 => (x"70",x"87",x"cc",x"e2"),
  2293 => (x"02",x"99",x"c2",x"49"),
  2294 => (x"c2",x"87",x"ed",x"c0"),
  2295 => (x"02",x"bf",x"ce",x"ec"),
  2296 => (x"c1",x"48",x"87",x"c9"),
  2297 => (x"d2",x"ec",x"c2",x"88"),
  2298 => (x"c2",x"87",x"d8",x"58"),
  2299 => (x"49",x"bf",x"ca",x"ec"),
  2300 => (x"66",x"c4",x"91",x"cc"),
  2301 => (x"7e",x"a1",x"c8",x"81"),
  2302 => (x"c0",x"02",x"bf",x"6e"),
  2303 => (x"ff",x"4b",x"87",x"c5"),
  2304 => (x"c8",x"0f",x"73",x"49"),
  2305 => (x"78",x"c1",x"48",x"a6"),
  2306 => (x"99",x"c4",x"49",x"74"),
  2307 => (x"c3",x"87",x"ce",x"05"),
  2308 => (x"ca",x"e1",x"49",x"f2"),
  2309 => (x"c2",x"49",x"70",x"87"),
  2310 => (x"fd",x"c0",x"02",x"99"),
  2311 => (x"48",x"a6",x"c8",x"87"),
  2312 => (x"bf",x"ca",x"ec",x"c2"),
  2313 => (x"49",x"66",x"c8",x"78"),
  2314 => (x"ec",x"c2",x"89",x"c1"),
  2315 => (x"6e",x"7e",x"bf",x"ce"),
  2316 => (x"c0",x"06",x"a9",x"b7"),
  2317 => (x"c1",x"48",x"87",x"c9"),
  2318 => (x"d2",x"ec",x"c2",x"80"),
  2319 => (x"c8",x"87",x"d6",x"58"),
  2320 => (x"91",x"cc",x"49",x"66"),
  2321 => (x"c8",x"81",x"66",x"c4"),
  2322 => (x"bf",x"6e",x"7e",x"a1"),
  2323 => (x"87",x"c5",x"c0",x"02"),
  2324 => (x"73",x"49",x"fe",x"4b"),
  2325 => (x"48",x"a6",x"c8",x"0f"),
  2326 => (x"fd",x"c3",x"78",x"c1"),
  2327 => (x"fe",x"df",x"ff",x"49"),
  2328 => (x"c2",x"49",x"70",x"87"),
  2329 => (x"ee",x"c0",x"02",x"99"),
  2330 => (x"ce",x"ec",x"c2",x"87"),
  2331 => (x"c9",x"c0",x"02",x"bf"),
  2332 => (x"ce",x"ec",x"c2",x"87"),
  2333 => (x"c0",x"78",x"c0",x"48"),
  2334 => (x"ec",x"c2",x"87",x"d8"),
  2335 => (x"cc",x"49",x"bf",x"ca"),
  2336 => (x"81",x"66",x"c4",x"91"),
  2337 => (x"6e",x"7e",x"a1",x"c8"),
  2338 => (x"c5",x"c0",x"02",x"bf"),
  2339 => (x"49",x"fd",x"4b",x"87"),
  2340 => (x"a6",x"c8",x"0f",x"73"),
  2341 => (x"c3",x"78",x"c1",x"48"),
  2342 => (x"df",x"ff",x"49",x"fa"),
  2343 => (x"49",x"70",x"87",x"c1"),
  2344 => (x"c1",x"02",x"99",x"c2"),
  2345 => (x"a6",x"c8",x"87",x"c0"),
  2346 => (x"ca",x"ec",x"c2",x"48"),
  2347 => (x"66",x"c8",x"78",x"bf"),
  2348 => (x"c4",x"88",x"c1",x"48"),
  2349 => (x"ec",x"c2",x"58",x"a6"),
  2350 => (x"6e",x"48",x"bf",x"ce"),
  2351 => (x"c0",x"03",x"a8",x"b7"),
  2352 => (x"ec",x"c2",x"87",x"c9"),
  2353 => (x"78",x"6e",x"48",x"ce"),
  2354 => (x"c8",x"87",x"d6",x"c0"),
  2355 => (x"91",x"cc",x"49",x"66"),
  2356 => (x"c8",x"81",x"66",x"c4"),
  2357 => (x"bf",x"6e",x"7e",x"a1"),
  2358 => (x"87",x"c5",x"c0",x"02"),
  2359 => (x"73",x"49",x"fc",x"4b"),
  2360 => (x"48",x"a6",x"c8",x"0f"),
  2361 => (x"ec",x"c2",x"78",x"c1"),
  2362 => (x"c0",x"4a",x"bf",x"ce"),
  2363 => (x"c0",x"06",x"aa",x"b7"),
  2364 => (x"8a",x"c1",x"87",x"c9"),
  2365 => (x"01",x"aa",x"b7",x"c0"),
  2366 => (x"74",x"87",x"f7",x"ff"),
  2367 => (x"99",x"f0",x"c3",x"49"),
  2368 => (x"87",x"cf",x"c0",x"05"),
  2369 => (x"ff",x"49",x"da",x"c1"),
  2370 => (x"70",x"87",x"d4",x"dd"),
  2371 => (x"02",x"99",x"c2",x"49"),
  2372 => (x"c2",x"87",x"ce",x"c1"),
  2373 => (x"7e",x"bf",x"c6",x"ec"),
  2374 => (x"c2",x"48",x"a6",x"c4"),
  2375 => (x"78",x"bf",x"ce",x"ec"),
  2376 => (x"48",x"4a",x"66",x"c4"),
  2377 => (x"06",x"a8",x"b7",x"c0"),
  2378 => (x"6e",x"87",x"d0",x"c0"),
  2379 => (x"c4",x"80",x"cc",x"48"),
  2380 => (x"8a",x"c1",x"58",x"a6"),
  2381 => (x"01",x"aa",x"b7",x"c0"),
  2382 => (x"6e",x"87",x"f0",x"ff"),
  2383 => (x"c2",x"4b",x"bf",x"97"),
  2384 => (x"d1",x"c0",x"02",x"8b"),
  2385 => (x"c0",x"05",x"8b",x"87"),
  2386 => (x"4a",x"6e",x"87",x"d7"),
  2387 => (x"49",x"6a",x"82",x"c8"),
  2388 => (x"c0",x"87",x"c2",x"f5"),
  2389 => (x"4b",x"6e",x"87",x"cb"),
  2390 => (x"4b",x"6b",x"83",x"c8"),
  2391 => (x"73",x"49",x"66",x"c4"),
  2392 => (x"02",x"9d",x"75",x"0f"),
  2393 => (x"6d",x"87",x"e9",x"c0"),
  2394 => (x"87",x"e4",x"c0",x"02"),
  2395 => (x"db",x"ff",x"49",x"6d"),
  2396 => (x"49",x"70",x"87",x"ed"),
  2397 => (x"c0",x"02",x"99",x"c1"),
  2398 => (x"a5",x"c4",x"87",x"cb"),
  2399 => (x"ce",x"ec",x"c2",x"4b"),
  2400 => (x"4b",x"6b",x"49",x"bf"),
  2401 => (x"02",x"85",x"c8",x"0f"),
  2402 => (x"6d",x"87",x"c5",x"c0"),
  2403 => (x"87",x"dc",x"ff",x"05"),
  2404 => (x"c0",x"02",x"66",x"c8"),
  2405 => (x"ec",x"c2",x"87",x"c8"),
  2406 => (x"f1",x"49",x"bf",x"ce"),
  2407 => (x"8e",x"f4",x"87",x"e0"),
  2408 => (x"58",x"87",x"ea",x"f3"),
  2409 => (x"1d",x"14",x"11",x"12"),
  2410 => (x"5a",x"23",x"1c",x"1b"),
  2411 => (x"f5",x"94",x"91",x"59"),
  2412 => (x"00",x"f4",x"eb",x"f2"),
  2413 => (x"00",x"00",x"00",x"00"),
  2414 => (x"00",x"00",x"00",x"00"),
  2415 => (x"58",x"00",x"00",x"00"),
  2416 => (x"1d",x"11",x"14",x"12"),
  2417 => (x"5a",x"23",x"1c",x"1b"),
  2418 => (x"f5",x"91",x"94",x"59"),
  2419 => (x"00",x"f4",x"eb",x"f2"),
  2420 => (x"00",x"00",x"25",x"d4"),
  2421 => (x"4f",x"54",x"55",x"41"),
  2422 => (x"54",x"4f",x"4f",x"42"),
  2423 => (x"00",x"53",x"45",x"4e"),
  2424 => (x"00",x"00",x"19",x"d4"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

