library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f8c6c387",
    12 => x"86c0d04e",
    13 => x"49f8c6c3",
    14 => x"48c8f2c2",
    15 => x"0389d089",
    16 => x"404040c0",
    17 => x"d087f640",
    18 => x"50c00581",
    19 => x"f90589c1",
    20 => x"c7f2c287",
    21 => x"c3f2c24d",
    22 => x"02ad744c",
    23 => x"0f2487c4",
    24 => x"f7c187f7",
    25 => x"f2c287fe",
    26 => x"f2c24dc7",
    27 => x"ad744cc7",
    28 => x"c487c602",
    29 => x"f50f6c8c",
    30 => x"87fd0087",
    31 => x"5c5b5e0e",
    32 => x"86f00e5d",
    33 => x"a6c44cc0",
    34 => x"c078c048",
    35 => x"c04ba6e4",
    36 => x"484966e0",
    37 => x"e4c080c1",
    38 => x"481158a6",
    39 => x"7058a6c4",
    40 => x"f6c30298",
    41 => x"0266c487",
    42 => x"c487c6c3",
    43 => x"78c048a6",
    44 => x"f0c04a6e",
    45 => x"dac2028a",
    46 => x"8af3c087",
    47 => x"87dbc202",
    48 => x"dc028ac1",
    49 => x"028ac887",
    50 => x"c487c8c2",
    51 => x"87d1028a",
    52 => x"c1028ac3",
    53 => x"8ac287eb",
    54 => x"c387c602",
    55 => x"c9c2058a",
    56 => x"7383c487",
    57 => x"6989c449",
    58 => x"c1026e7e",
    59 => x"a6c887c8",
    60 => x"c478c048",
    61 => x"cc78c080",
    62 => x"4a6e4d66",
    63 => x"cf2ab7dc",
    64 => x"c4486e9a",
    65 => x"7258a630",
    66 => x"87c5029a",
    67 => x"c148a6c8",
    68 => x"06aac978",
    69 => x"f7c087c5",
    70 => x"c087c382",
    71 => x"66c882f0",
    72 => x"7287c702",
    73 => x"87f3c249",
    74 => x"85c184c1",
    75 => x"04adb7c8",
    76 => x"c187c7ff",
    77 => x"f0c087cf",
    78 => x"87dfc249",
    79 => x"c4c184c1",
    80 => x"7383c487",
    81 => x"6a8ac44a",
    82 => x"87dbc149",
    83 => x"4ca44970",
    84 => x"c487f2c0",
    85 => x"78c148a6",
    86 => x"c487eac0",
    87 => x"c44a7383",
    88 => x"c1496a8a",
    89 => x"84c187f5",
    90 => x"496e87db",
    91 => x"d487ecc1",
    92 => x"c0486e87",
    93 => x"c705a8e5",
    94 => x"48a6c487",
    95 => x"87c578c1",
    96 => x"d6c1496e",
    97 => x"66e0c087",
    98 => x"80c14849",
    99 => x"58a6e4c0",
   100 => x"a6c44811",
   101 => x"05987058",
   102 => x"7487cafc",
   103 => x"268ef048",
   104 => x"264c264d",
   105 => x"0e4f264b",
   106 => x"0e5c5b5e",
   107 => x"4cc04b71",
   108 => x"029a4a13",
   109 => x"497287cd",
   110 => x"c187e0c0",
   111 => x"9a4a1384",
   112 => x"7487f305",
   113 => x"264c2648",
   114 => x"1e4f264b",
   115 => x"73814873",
   116 => x"87c502a9",
   117 => x"f6055312",
   118 => x"1e4f2687",
   119 => x"4ac0ff1e",
   120 => x"c0c4486a",
   121 => x"58a6c498",
   122 => x"f3029870",
   123 => x"487a7187",
   124 => x"1e4f2626",
   125 => x"d4ff1e73",
   126 => x"7bffc34b",
   127 => x"ffc34a6b",
   128 => x"c8496b7b",
   129 => x"c3b17232",
   130 => x"4a6b7bff",
   131 => x"b27131c8",
   132 => x"6b7bffc3",
   133 => x"7232c849",
   134 => x"c44871b1",
   135 => x"264d2687",
   136 => x"264b264c",
   137 => x"5b5e0e4f",
   138 => x"710e5d5c",
   139 => x"4cd4ff4a",
   140 => x"ffc34872",
   141 => x"c27c7098",
   142 => x"05bfc8f2",
   143 => x"66d087c8",
   144 => x"d430c948",
   145 => x"66d058a6",
   146 => x"7129d849",
   147 => x"98ffc348",
   148 => x"66d07c70",
   149 => x"7129d049",
   150 => x"98ffc348",
   151 => x"66d07c70",
   152 => x"7129c849",
   153 => x"98ffc348",
   154 => x"66d07c70",
   155 => x"98ffc348",
   156 => x"49727c70",
   157 => x"487129d0",
   158 => x"7098ffc3",
   159 => x"c94b6c7c",
   160 => x"c34dfff0",
   161 => x"d005abff",
   162 => x"7cffc387",
   163 => x"8dc14b6c",
   164 => x"c387c602",
   165 => x"f002abff",
   166 => x"fd487387",
   167 => x"c01e87ff",
   168 => x"48d4ff49",
   169 => x"c178ffc3",
   170 => x"b7c8c381",
   171 => x"87f104a9",
   172 => x"731e4f26",
   173 => x"c487e71e",
   174 => x"c04bdff8",
   175 => x"f0ffc01e",
   176 => x"fd49f7c1",
   177 => x"86c487df",
   178 => x"c005a8c1",
   179 => x"d4ff87ea",
   180 => x"78ffc348",
   181 => x"c0c0c0c1",
   182 => x"c01ec0c0",
   183 => x"e9c1f0e1",
   184 => x"87c1fd49",
   185 => x"987086c4",
   186 => x"ff87ca05",
   187 => x"ffc348d4",
   188 => x"cb48c178",
   189 => x"87e6fe87",
   190 => x"fe058bc1",
   191 => x"48c087fd",
   192 => x"1e87defc",
   193 => x"d4ff1e73",
   194 => x"78ffc348",
   195 => x"fa49fecc",
   196 => x"4bd387d5",
   197 => x"ffc01ec0",
   198 => x"49c1c1f0",
   199 => x"c487c6fc",
   200 => x"05987086",
   201 => x"d4ff87ca",
   202 => x"78ffc348",
   203 => x"87cb48c1",
   204 => x"c187ebfd",
   205 => x"dbff058b",
   206 => x"fb48c087",
   207 => x"4d4387e3",
   208 => x"4d430044",
   209 => x"20383544",
   210 => x"200a6425",
   211 => x"4d430020",
   212 => x"5f383544",
   213 => x"64252032",
   214 => x"0020200a",
   215 => x"35444d43",
   216 => x"64252038",
   217 => x"0020200a",
   218 => x"43484453",
   219 => x"696e4920",
   220 => x"6c616974",
   221 => x"74617a69",
   222 => x"206e6f69",
   223 => x"6f727265",
   224 => x"000a2172",
   225 => x"5f646d63",
   226 => x"38444d43",
   227 => x"73657220",
   228 => x"736e6f70",
   229 => x"25203a65",
   230 => x"49000a64",
   231 => x"00525245",
   232 => x"00495053",
   233 => x"63204453",
   234 => x"20647261",
   235 => x"657a6973",
   236 => x"20736920",
   237 => x"000a6425",
   238 => x"74697257",
   239 => x"61662065",
   240 => x"64656c69",
   241 => x"5f63000a",
   242 => x"657a6973",
   243 => x"6c756d5f",
   244 => x"25203a74",
   245 => x"72202c64",
   246 => x"5f646165",
   247 => x"6c5f6c62",
   248 => x"203a6e65",
   249 => x"202c6425",
   250 => x"7a697363",
   251 => x"25203a65",
   252 => x"4d000a64",
   253 => x"20746c75",
   254 => x"000a6425",
   255 => x"62206425",
   256 => x"6b636f6c",
   257 => x"666f2073",
   258 => x"7a697320",
   259 => x"64252065",
   260 => x"6425000a",
   261 => x"6f6c6220",
   262 => x"20736b63",
   263 => x"3520666f",
   264 => x"62203231",
   265 => x"73657479",
   266 => x"5e0e000a",
   267 => x"0e5d5c5b",
   268 => x"f94dd4ff",
   269 => x"eac687e8",
   270 => x"f0e1c01e",
   271 => x"f749c8c1",
   272 => x"4b7087e3",
   273 => x"1ec4ce1e",
   274 => x"cc87f1f0",
   275 => x"02abc186",
   276 => x"eefa87c8",
   277 => x"c248c087",
   278 => x"d6f687ca",
   279 => x"cf497087",
   280 => x"c699ffff",
   281 => x"c802a9ea",
   282 => x"87d7fa87",
   283 => x"f3c148c0",
   284 => x"7dffc387",
   285 => x"f84cf1c0",
   286 => x"987087f8",
   287 => x"87cbc102",
   288 => x"ffc01ec0",
   289 => x"49fac1f0",
   290 => x"c487daf6",
   291 => x"9b4b7086",
   292 => x"87edc005",
   293 => x"1ec2cd1e",
   294 => x"c387e1ef",
   295 => x"4b6d7dff",
   296 => x"1ececd1e",
   297 => x"d087d5ef",
   298 => x"7dffc386",
   299 => x"737d7d7d",
   300 => x"99c0c149",
   301 => x"c187c502",
   302 => x"87e8c048",
   303 => x"e3c048c0",
   304 => x"cd1e7387",
   305 => x"f3ee1edc",
   306 => x"c286c887",
   307 => x"87cc05ac",
   308 => x"ee1ee8cd",
   309 => x"86c487e6",
   310 => x"87c848c0",
   311 => x"fe058cc1",
   312 => x"48c087d5",
   313 => x"0e87f6f4",
   314 => x"5d5c5b5e",
   315 => x"d0ff1e0e",
   316 => x"c0c0c84d",
   317 => x"c8f2c24b",
   318 => x"ce78c148",
   319 => x"e6f249e0",
   320 => x"6d4cc787",
   321 => x"c4987348",
   322 => x"987058a6",
   323 => x"6d87cc02",
   324 => x"c4987348",
   325 => x"987058a6",
   326 => x"c287f405",
   327 => x"87fef57d",
   328 => x"9873486d",
   329 => x"7058a6c4",
   330 => x"87cc0298",
   331 => x"9873486d",
   332 => x"7058a6c4",
   333 => x"87f40598",
   334 => x"1ec07dc3",
   335 => x"c1d0e5c0",
   336 => x"e0f349c0",
   337 => x"c186c487",
   338 => x"87c105a8",
   339 => x"05acc24c",
   340 => x"dbce87cb",
   341 => x"87cff149",
   342 => x"d8c148c0",
   343 => x"058cc187",
   344 => x"fb87e0fe",
   345 => x"f2c287c4",
   346 => x"987058cc",
   347 => x"c187cd05",
   348 => x"f0ffc01e",
   349 => x"f249d0c1",
   350 => x"86c487eb",
   351 => x"c348d4ff",
   352 => x"e7c578ff",
   353 => x"d0f2c287",
   354 => x"ce1e7058",
   355 => x"ebeb1ee4",
   356 => x"6d86c887",
   357 => x"c4987348",
   358 => x"987058a6",
   359 => x"6d87cc02",
   360 => x"c4987348",
   361 => x"987058a6",
   362 => x"c287f405",
   363 => x"48d4ff7d",
   364 => x"c178ffc3",
   365 => x"e4f12648",
   366 => x"5b5e0e87",
   367 => x"1e0e5d5c",
   368 => x"4bc0c0c8",
   369 => x"eec54cc0",
   370 => x"c44adfcd",
   371 => x"d4ff5ca6",
   372 => x"7cffc34c",
   373 => x"fec3486c",
   374 => x"c0c205a8",
   375 => x"05997187",
   376 => x"ff87e2c0",
   377 => x"7348bfd0",
   378 => x"58a6c498",
   379 => x"ce029870",
   380 => x"bfd0ff87",
   381 => x"c4987348",
   382 => x"987058a6",
   383 => x"ff87f205",
   384 => x"d1c448d0",
   385 => x"4866d478",
   386 => x"06a8b7c0",
   387 => x"c387e0c0",
   388 => x"4a6c7cff",
   389 => x"c7029971",
   390 => x"970a7187",
   391 => x"81c10a7a",
   392 => x"c14866d4",
   393 => x"58a6d888",
   394 => x"01a8b7c0",
   395 => x"c387e0ff",
   396 => x"717c7cff",
   397 => x"e1c00599",
   398 => x"bfd0ff87",
   399 => x"c4987348",
   400 => x"987058a6",
   401 => x"ff87ce02",
   402 => x"7348bfd0",
   403 => x"58a6c498",
   404 => x"f2059870",
   405 => x"48d0ff87",
   406 => x"4ac178d0",
   407 => x"058ac17e",
   408 => x"6e87eefd",
   409 => x"f4ee2648",
   410 => x"5b5e0e87",
   411 => x"711e0e5c",
   412 => x"c0c0c84a",
   413 => x"ff4cc04b",
   414 => x"ffc348d4",
   415 => x"bfd0ff78",
   416 => x"c4987348",
   417 => x"987058a6",
   418 => x"ff87ce02",
   419 => x"7348bfd0",
   420 => x"58a6c498",
   421 => x"f2059870",
   422 => x"48d0ff87",
   423 => x"ff78c3c4",
   424 => x"ffc348d4",
   425 => x"c01e7278",
   426 => x"d1c1f0ff",
   427 => x"87f5ed49",
   428 => x"987086c4",
   429 => x"87eec005",
   430 => x"d41ec0c8",
   431 => x"f8fb4966",
   432 => x"7086c487",
   433 => x"bfd0ff4c",
   434 => x"c4987348",
   435 => x"987058a6",
   436 => x"ff87ce02",
   437 => x"7348bfd0",
   438 => x"58a6c498",
   439 => x"f2059870",
   440 => x"48d0ff87",
   441 => x"487478c2",
   442 => x"87f3ec26",
   443 => x"5c5b5e0e",
   444 => x"c01e0e5d",
   445 => x"f0ffc01e",
   446 => x"ec49c9c1",
   447 => x"1ed287e7",
   448 => x"49d6f2c2",
   449 => x"c887f2fa",
   450 => x"c14dc086",
   451 => x"adb7d285",
   452 => x"c287f804",
   453 => x"bf97d6f2",
   454 => x"99c0c349",
   455 => x"05a9c0c1",
   456 => x"c287e7c0",
   457 => x"bf97ddf2",
   458 => x"c231d049",
   459 => x"bf97def2",
   460 => x"7232c84a",
   461 => x"dff2c2b1",
   462 => x"b14abf97",
   463 => x"ffcf4d71",
   464 => x"c19dffff",
   465 => x"c235ca85",
   466 => x"f2c287de",
   467 => x"4bbf97df",
   468 => x"9bc633c1",
   469 => x"97e0f2c2",
   470 => x"b7c749bf",
   471 => x"c2b37129",
   472 => x"bf97dbf2",
   473 => x"98cf4849",
   474 => x"c258a6c4",
   475 => x"bf97dcf2",
   476 => x"ca9cc34c",
   477 => x"ddf2c234",
   478 => x"c249bf97",
   479 => x"c2b47131",
   480 => x"bf97def2",
   481 => x"99c0c349",
   482 => x"7129b7c6",
   483 => x"701e74b4",
   484 => x"cf1e731e",
   485 => x"e3e31ec6",
   486 => x"c183c287",
   487 => x"70307348",
   488 => x"f3cf1e4b",
   489 => x"87d4e31e",
   490 => x"66d848c1",
   491 => x"58a6dc30",
   492 => x"4d49a4c1",
   493 => x"1e709573",
   494 => x"fccf1e75",
   495 => x"87fce21e",
   496 => x"6e86e4c0",
   497 => x"b7c0c848",
   498 => x"87d206a8",
   499 => x"486e35c1",
   500 => x"c428b7c1",
   501 => x"c0c858a6",
   502 => x"ff01a8b7",
   503 => x"1e7587ee",
   504 => x"e21ed2d0",
   505 => x"86c887d6",
   506 => x"e8264875",
   507 => x"5e0e87ef",
   508 => x"710e5c5b",
   509 => x"d04cc04b",
   510 => x"b7c04866",
   511 => x"e3c006a8",
   512 => x"cc4a1387",
   513 => x"49bf9766",
   514 => x"c14866cc",
   515 => x"58a6d080",
   516 => x"02aab771",
   517 => x"48c187c4",
   518 => x"84c187cc",
   519 => x"acb766d0",
   520 => x"87ddff04",
   521 => x"87c248c0",
   522 => x"4c264d26",
   523 => x"4f264b26",
   524 => x"5c5b5e0e",
   525 => x"fac20e5d",
   526 => x"78c048fc",
   527 => x"49ddefc0",
   528 => x"c287e4e5",
   529 => x"c01ef4f2",
   530 => x"87ddf849",
   531 => x"987086c4",
   532 => x"c087cc05",
   533 => x"e549c9ec",
   534 => x"48c087cd",
   535 => x"c087e7ca",
   536 => x"e549eaef",
   537 => x"4bc087c1",
   538 => x"48f4ffc2",
   539 => x"1ec878c1",
   540 => x"1ec1f0c0",
   541 => x"49eaf3c2",
   542 => x"c887f3fd",
   543 => x"05987086",
   544 => x"ffc287c6",
   545 => x"78c048f4",
   546 => x"f0c01ec8",
   547 => x"f4c21eca",
   548 => x"d9fd49c6",
   549 => x"7086c887",
   550 => x"87c60598",
   551 => x"48f4ffc2",
   552 => x"ffc278c0",
   553 => x"c01ebff4",
   554 => x"ff1ed3f0",
   555 => x"c887cddf",
   556 => x"f4ffc286",
   557 => x"f7c102bf",
   558 => x"f2fac287",
   559 => x"1e49bf9f",
   560 => x"49f2fac2",
   561 => x"a0c2f848",
   562 => x"d01e7189",
   563 => x"1ec0c81e",
   564 => x"1efbecc0",
   565 => x"87e4deff",
   566 => x"f9c286d4",
   567 => x"c24bbffa",
   568 => x"bf9ff2fa",
   569 => x"ead6c54a",
   570 => x"c8c005aa",
   571 => x"faf9c287",
   572 => x"d4c04bbf",
   573 => x"d5e9ca87",
   574 => x"ccc002aa",
   575 => x"ddecc087",
   576 => x"87e3e249",
   577 => x"fdc748c0",
   578 => x"c01e7387",
   579 => x"ff1ef8ed",
   580 => x"c287e9dd",
   581 => x"731ef4f2",
   582 => x"87cdf549",
   583 => x"987086cc",
   584 => x"87c5c005",
   585 => x"ddc748c0",
   586 => x"d0eec087",
   587 => x"87f7e149",
   588 => x"1ee6f0c0",
   589 => x"87c4ddff",
   590 => x"f0c01ec8",
   591 => x"f4c21efe",
   592 => x"e9fa49c6",
   593 => x"7086cc87",
   594 => x"c9c00598",
   595 => x"fcfac287",
   596 => x"c078c148",
   597 => x"1ec887e4",
   598 => x"1ec7f1c0",
   599 => x"49eaf3c2",
   600 => x"c887cbfa",
   601 => x"02987086",
   602 => x"c087cfc0",
   603 => x"ff1ef7ee",
   604 => x"c487c9dc",
   605 => x"c648c086",
   606 => x"fac287cc",
   607 => x"49bf97f2",
   608 => x"05a9d5c1",
   609 => x"c287cdc0",
   610 => x"bf97f3fa",
   611 => x"a9eac249",
   612 => x"87c5c002",
   613 => x"edc548c0",
   614 => x"f4f2c287",
   615 => x"c34cbf97",
   616 => x"c002ace9",
   617 => x"ebc387cc",
   618 => x"c5c002ac",
   619 => x"c548c087",
   620 => x"f2c287d4",
   621 => x"49bf97ff",
   622 => x"ccc00599",
   623 => x"c0f3c287",
   624 => x"c249bf97",
   625 => x"c5c002a9",
   626 => x"c448c087",
   627 => x"f3c287f8",
   628 => x"48bf97c1",
   629 => x"58f8fac2",
   630 => x"c14a4970",
   631 => x"fcfac28a",
   632 => x"711e725a",
   633 => x"d0f1c01e",
   634 => x"cfdaff1e",
   635 => x"c286cc87",
   636 => x"bf97c2f3",
   637 => x"c2817349",
   638 => x"bf97c3f3",
   639 => x"35c84d4a",
   640 => x"ffc28571",
   641 => x"f3c25dd4",
   642 => x"48bf97c4",
   643 => x"58e8ffc2",
   644 => x"bffcfac2",
   645 => x"87dcc202",
   646 => x"efc01ec8",
   647 => x"f4c21ed4",
   648 => x"c9f749c6",
   649 => x"7086c887",
   650 => x"c5c00298",
   651 => x"c348c087",
   652 => x"fac287d4",
   653 => x"484abff4",
   654 => x"fbc230c4",
   655 => x"ffc258c4",
   656 => x"f3c25ae4",
   657 => x"49bf97d9",
   658 => x"f3c231c8",
   659 => x"4bbf97d8",
   660 => x"f3c249a1",
   661 => x"4bbf97da",
   662 => x"a17333d0",
   663 => x"dbf3c249",
   664 => x"d84bbf97",
   665 => x"49a17333",
   666 => x"59ecffc2",
   667 => x"bfe4ffc2",
   668 => x"d0ffc291",
   669 => x"ffc281bf",
   670 => x"f3c259d8",
   671 => x"4bbf97e1",
   672 => x"f3c233c8",
   673 => x"4cbf97e0",
   674 => x"f3c24ba3",
   675 => x"4cbf97e2",
   676 => x"a37434d0",
   677 => x"e3f3c24b",
   678 => x"cf4cbf97",
   679 => x"7434d89c",
   680 => x"ffc24ba3",
   681 => x"8bc25bdc",
   682 => x"ffc29273",
   683 => x"a17248dc",
   684 => x"87cbc178",
   685 => x"97c6f3c2",
   686 => x"31c849bf",
   687 => x"97c5f3c2",
   688 => x"49a14abf",
   689 => x"59c4fbc2",
   690 => x"ffc731c5",
   691 => x"c229c981",
   692 => x"c259e4ff",
   693 => x"bf97cbf3",
   694 => x"c232c84a",
   695 => x"bf97caf3",
   696 => x"c24aa24b",
   697 => x"c25aecff",
   698 => x"92bfe4ff",
   699 => x"ffc28275",
   700 => x"ffc25ae0",
   701 => x"78c048d8",
   702 => x"48d4ffc2",
   703 => x"c078a172",
   704 => x"87e3cd49",
   705 => x"dff448c1",
   706 => x"61655287",
   707 => x"666f2064",
   708 => x"52424d20",
   709 => x"69616620",
   710 => x"0a64656c",
   711 => x"206f4e00",
   712 => x"74726170",
   713 => x"6f697469",
   714 => x"6973206e",
   715 => x"74616e67",
   716 => x"20657275",
   717 => x"6e756f66",
   718 => x"4d000a64",
   719 => x"69735242",
   720 => x"203a657a",
   721 => x"202c6425",
   722 => x"74726170",
   723 => x"6f697469",
   724 => x"7a69736e",
   725 => x"25203a65",
   726 => x"6f202c64",
   727 => x"65736666",
   728 => x"666f2074",
   729 => x"67697320",
   730 => x"6425203a",
   731 => x"6973202c",
   732 => x"78302067",
   733 => x"000a7825",
   734 => x"64616552",
   735 => x"20676e69",
   736 => x"746f6f62",
   737 => x"63657320",
   738 => x"20726f74",
   739 => x"000a6425",
   740 => x"64616552",
   741 => x"6f6f6220",
   742 => x"65732074",
   743 => x"726f7463",
   744 => x"6f726620",
   745 => x"6966206d",
   746 => x"20747372",
   747 => x"74726170",
   748 => x"6f697469",
   749 => x"55000a6e",
   750 => x"7075736e",
   751 => x"74726f70",
   752 => x"70206465",
   753 => x"69747261",
   754 => x"6e6f6974",
   755 => x"70797420",
   756 => x"000d2165",
   757 => x"33544146",
   758 => x"20202032",
   759 => x"61655200",
   760 => x"676e6964",
   761 => x"52424d20",
   762 => x"424d000a",
   763 => x"75732052",
   764 => x"73656363",
   765 => x"6c756673",
   766 => x"7220796c",
   767 => x"0a646165",
   768 => x"54414600",
   769 => x"20203631",
   770 => x"41460020",
   771 => x"20323354",
   772 => x"50002020",
   773 => x"69747261",
   774 => x"6e6f6974",
   775 => x"6e756f63",
   776 => x"64252074",
   777 => x"7548000a",
   778 => x"6e69746e",
   779 => x"6f662067",
   780 => x"69662072",
   781 => x"7973656c",
   782 => x"6d657473",
   783 => x"4146000a",
   784 => x"20323354",
   785 => x"46002020",
   786 => x"36315441",
   787 => x"00202020",
   788 => x"73756c43",
   789 => x"20726574",
   790 => x"657a6973",
   791 => x"6425203a",
   792 => x"6c43202c",
   793 => x"65747375",
   794 => x"616d2072",
   795 => x"202c6b73",
   796 => x"000a6425",
   797 => x"6e65704f",
   798 => x"66206465",
   799 => x"2c656c69",
   800 => x"616f6c20",
   801 => x"676e6964",
   802 => x"0a2e2e2e",
   803 => x"6e614300",
   804 => x"6f207427",
   805 => x"206e6570",
   806 => x"000a7325",
   807 => x"5c5b5e0e",
   808 => x"4a710e5d",
   809 => x"bffcfac2",
   810 => x"7287cc02",
   811 => x"2bb7c74b",
   812 => x"ffc14d72",
   813 => x"7287ca9d",
   814 => x"2bb7c84b",
   815 => x"ffc34d72",
   816 => x"f4f2c29d",
   817 => x"d0ffc21e",
   818 => x"817349bf",
   819 => x"87d9e671",
   820 => x"987086c4",
   821 => x"c087c505",
   822 => x"87e6c048",
   823 => x"bffcfac2",
   824 => x"7587d202",
   825 => x"c291c449",
   826 => x"6981f4f2",
   827 => x"ffffcf4c",
   828 => x"cb9cffff",
   829 => x"c2497587",
   830 => x"f4f2c291",
   831 => x"4c699f81",
   832 => x"e3ec4874",
   833 => x"5b5e0e87",
   834 => x"f40e5d5c",
   835 => x"c04c7186",
   836 => x"ecffc24b",
   837 => x"a6c47ebf",
   838 => x"f0ffc248",
   839 => x"a6c878bf",
   840 => x"c278c048",
   841 => x"48bfc0fb",
   842 => x"c206a8c0",
   843 => x"66c887e3",
   844 => x"0599cf49",
   845 => x"f2c287d8",
   846 => x"66c81ef4",
   847 => x"80c14849",
   848 => x"e458a6cc",
   849 => x"86c487e3",
   850 => x"4bf4f2c2",
   851 => x"e0c087c3",
   852 => x"4a6b9783",
   853 => x"e7c1029a",
   854 => x"aae5c387",
   855 => x"87e0c102",
   856 => x"9749a3cb",
   857 => x"99d84969",
   858 => x"87d4c105",
   859 => x"d0ff4973",
   860 => x"1ecb87f5",
   861 => x"1e66e0c0",
   862 => x"f1e94973",
   863 => x"7086c887",
   864 => x"fbc00598",
   865 => x"4aa3dc87",
   866 => x"6a49a4c4",
   867 => x"49a3da79",
   868 => x"9f4da4c8",
   869 => x"c27d4869",
   870 => x"02bffcfa",
   871 => x"a3d487d3",
   872 => x"49699f49",
   873 => x"99ffffc0",
   874 => x"30d04871",
   875 => x"c258a6c4",
   876 => x"6e7ec087",
   877 => x"70806d48",
   878 => x"c17cc07d",
   879 => x"87c5c148",
   880 => x"c14866c8",
   881 => x"58a6cc80",
   882 => x"bfc0fbc2",
   883 => x"ddfd04a8",
   884 => x"fcfac287",
   885 => x"eac002bf",
   886 => x"fa496e87",
   887 => x"a6c487fe",
   888 => x"cf497058",
   889 => x"f8ffffff",
   890 => x"d602a999",
   891 => x"c2497087",
   892 => x"f4fac289",
   893 => x"ffc291bf",
   894 => x"7148bfd4",
   895 => x"58a6c880",
   896 => x"c087dbfc",
   897 => x"e88ef448",
   898 => x"731e87de",
   899 => x"6a4a711e",
   900 => x"7181c149",
   901 => x"f8fac27a",
   902 => x"cb0599bf",
   903 => x"4ba2c887",
   904 => x"f7f9496b",
   905 => x"7b497087",
   906 => x"ffe748c1",
   907 => x"1e731e87",
   908 => x"ffc24b71",
   909 => x"c849bfd4",
   910 => x"4a6a4aa3",
   911 => x"fac28ac2",
   912 => x"7292bff4",
   913 => x"fac249a1",
   914 => x"6b4abff8",
   915 => x"49a1729a",
   916 => x"711e66c8",
   917 => x"c487d2e0",
   918 => x"05987086",
   919 => x"48c087c4",
   920 => x"48c187c2",
   921 => x"0e87c5e7",
   922 => x"0e5c5b5e",
   923 => x"4bc04a71",
   924 => x"c0029a72",
   925 => x"a2da87e0",
   926 => x"4b699f49",
   927 => x"bffcfac2",
   928 => x"d487cf02",
   929 => x"699f49a2",
   930 => x"ffc04c49",
   931 => x"34d09cff",
   932 => x"4cc087c2",
   933 => x"9b73b374",
   934 => x"4a87df02",
   935 => x"fac28ac2",
   936 => x"9249bff4",
   937 => x"bfd4ffc2",
   938 => x"c2807248",
   939 => x"7158f4ff",
   940 => x"c230c448",
   941 => x"c058c4fb",
   942 => x"ffc287e9",
   943 => x"c24bbfd8",
   944 => x"c248f0ff",
   945 => x"78bfdcff",
   946 => x"bffcfac2",
   947 => x"c287c902",
   948 => x"49bff4fa",
   949 => x"87c731c4",
   950 => x"bfe0ffc2",
   951 => x"c231c449",
   952 => x"c259c4fb",
   953 => x"e55bf0ff",
   954 => x"5e0e87c0",
   955 => x"0e5d5c5b",
   956 => x"9a4a711e",
   957 => x"c287de02",
   958 => x"c048f0f2",
   959 => x"e8f2c278",
   960 => x"f0ffc248",
   961 => x"f2c278bf",
   962 => x"ffc248ec",
   963 => x"c178bfec",
   964 => x"c048e2c2",
   965 => x"c0fbc278",
   966 => x"f2c249bf",
   967 => x"714abff0",
   968 => x"fec303aa",
   969 => x"cf497287",
   970 => x"e1c00599",
   971 => x"f4f2c287",
   972 => x"e8f2c21e",
   973 => x"f2c249bf",
   974 => x"a1c148e8",
   975 => x"dcff7178",
   976 => x"86c487e7",
   977 => x"48dec2c1",
   978 => x"78f4f2c2",
   979 => x"c2c187cc",
   980 => x"c048bfde",
   981 => x"c2c180e0",
   982 => x"f2c258e2",
   983 => x"c148bff0",
   984 => x"f4f2c280",
   985 => x"dec2c158",
   986 => x"a3cb4bbf",
   987 => x"cf4c1149",
   988 => x"ddc105ac",
   989 => x"109e2787",
   990 => x"97bf0000",
   991 => x"99df49bf",
   992 => x"91cd89c1",
   993 => x"81c4fbc2",
   994 => x"124aa3c1",
   995 => x"4aa3c351",
   996 => x"a3c55112",
   997 => x"c751124a",
   998 => x"51124aa3",
   999 => x"124aa3c9",
  1000 => x"4aa3ce51",
  1001 => x"a3d05112",
  1002 => x"d251124a",
  1003 => x"51124aa3",
  1004 => x"124aa3d4",
  1005 => x"4aa3d651",
  1006 => x"a3d85112",
  1007 => x"dc51124a",
  1008 => x"51124aa3",
  1009 => x"124aa3de",
  1010 => x"e2c2c151",
  1011 => x"c178c148",
  1012 => x"497487c1",
  1013 => x"c00599c8",
  1014 => x"497487f3",
  1015 => x"d00599d0",
  1016 => x"0266d487",
  1017 => x"7387cac0",
  1018 => x"0f66d449",
  1019 => x"dc029870",
  1020 => x"e2c2c187",
  1021 => x"c6c005bf",
  1022 => x"c4fbc287",
  1023 => x"c150c048",
  1024 => x"c048e2c2",
  1025 => x"dec2c178",
  1026 => x"ccc248bf",
  1027 => x"e2c2c187",
  1028 => x"c278c048",
  1029 => x"49bfc0fb",
  1030 => x"bff0f2c2",
  1031 => x"04aa714a",
  1032 => x"c287c2fc",
  1033 => x"05bff0ff",
  1034 => x"c287c8c0",
  1035 => x"02bffcfa",
  1036 => x"c287e4c1",
  1037 => x"49bfecf2",
  1038 => x"c287e1f1",
  1039 => x"7058f0f2",
  1040 => x"fcfac24d",
  1041 => x"d7c002bf",
  1042 => x"cf497587",
  1043 => x"f8ffffff",
  1044 => x"c002a999",
  1045 => x"4cc087c5",
  1046 => x"c187d9c0",
  1047 => x"87d4c04c",
  1048 => x"ffcf4975",
  1049 => x"02a999f8",
  1050 => x"c087c5c0",
  1051 => x"87c2c07e",
  1052 => x"4c6e7ec1",
  1053 => x"c0059c74",
  1054 => x"497587dd",
  1055 => x"fac289c2",
  1056 => x"c291bff4",
  1057 => x"48bfd4ff",
  1058 => x"f2c28071",
  1059 => x"f2c258ec",
  1060 => x"78c048f0",
  1061 => x"c087fef9",
  1062 => x"deff2648",
  1063 => x"000087ca",
  1064 => x"00000000",
  1065 => x"ff1e0000",
  1066 => x"ffc348d4",
  1067 => x"99496878",
  1068 => x"c087c602",
  1069 => x"ee05a9fb",
  1070 => x"26487187",
  1071 => x"5b5e0e4f",
  1072 => x"4a710e5c",
  1073 => x"d4ff4bc0",
  1074 => x"78ffc348",
  1075 => x"02994968",
  1076 => x"c087c1c1",
  1077 => x"c002a9ec",
  1078 => x"fbc087fa",
  1079 => x"f3c002a9",
  1080 => x"b766cc87",
  1081 => x"87cc03ab",
  1082 => x"c70266d0",
  1083 => x"97097287",
  1084 => x"82c10979",
  1085 => x"c2029971",
  1086 => x"ff83c187",
  1087 => x"ffc348d4",
  1088 => x"99496878",
  1089 => x"c087cd02",
  1090 => x"c702a9ec",
  1091 => x"a9fbc087",
  1092 => x"87cdff05",
  1093 => x"c30266d0",
  1094 => x"7a97c087",
  1095 => x"05a9fbc0",
  1096 => x"4c7387c7",
  1097 => x"c28c0cc0",
  1098 => x"744c7387",
  1099 => x"2687c248",
  1100 => x"264c264d",
  1101 => x"1e4f264b",
  1102 => x"c348d4ff",
  1103 => x"496878ff",
  1104 => x"a9b7f0c0",
  1105 => x"c087ca04",
  1106 => x"01a9b7f9",
  1107 => x"f0c087c3",
  1108 => x"b7c1c189",
  1109 => x"87ca04a9",
  1110 => x"a9b7c6c1",
  1111 => x"c087c301",
  1112 => x"487189f7",
  1113 => x"5e0e4f26",
  1114 => x"0e5d5c5b",
  1115 => x"4c7186f4",
  1116 => x"c04bd4ff",
  1117 => x"ffc37e4d",
  1118 => x"bfd0ff7b",
  1119 => x"c0c0c848",
  1120 => x"58a6c898",
  1121 => x"d0029870",
  1122 => x"bfd0ff87",
  1123 => x"c0c0c848",
  1124 => x"58a6c898",
  1125 => x"f0059870",
  1126 => x"48d0ff87",
  1127 => x"d478e1c0",
  1128 => x"87c2fc7b",
  1129 => x"02994970",
  1130 => x"c387c7c1",
  1131 => x"a6c87bff",
  1132 => x"c8786b48",
  1133 => x"fbc04866",
  1134 => x"87c802a8",
  1135 => x"bfccc0c3",
  1136 => x"87eec002",
  1137 => x"99714dc1",
  1138 => x"87e6c002",
  1139 => x"02a9fbc0",
  1140 => x"d1fb87c3",
  1141 => x"7bffc387",
  1142 => x"c6c1496b",
  1143 => x"87cc05a9",
  1144 => x"7b7bffc3",
  1145 => x"6b48a6c8",
  1146 => x"4d49c078",
  1147 => x"ff059971",
  1148 => x"9d7587da",
  1149 => x"87dec105",
  1150 => x"6b7bffc3",
  1151 => x"7bffc34a",
  1152 => x"6b48a6c4",
  1153 => x"c1486e78",
  1154 => x"58a6c480",
  1155 => x"9749a4c8",
  1156 => x"66c84969",
  1157 => x"87da05a9",
  1158 => x"9749a4c9",
  1159 => x"05aa4969",
  1160 => x"a4ca87d0",
  1161 => x"49699749",
  1162 => x"05a966c4",
  1163 => x"4dc187c4",
  1164 => x"66c887d6",
  1165 => x"a8ecc048",
  1166 => x"c887c902",
  1167 => x"fbc04866",
  1168 => x"87c405a8",
  1169 => x"4dc17ec0",
  1170 => x"c87bffc3",
  1171 => x"786b48a6",
  1172 => x"fe029d75",
  1173 => x"d0ff87e2",
  1174 => x"c0c848bf",
  1175 => x"a6c898c0",
  1176 => x"02987058",
  1177 => x"d0ff87d0",
  1178 => x"c0c848bf",
  1179 => x"a6c898c0",
  1180 => x"05987058",
  1181 => x"d0ff87f0",
  1182 => x"78e0c048",
  1183 => x"8ef4486e",
  1184 => x"0e87ecfa",
  1185 => x"5d5c5b5e",
  1186 => x"d0ff1e0e",
  1187 => x"c0c0c84b",
  1188 => x"d4c0c34a",
  1189 => x"486b4dbf",
  1190 => x"a6c49872",
  1191 => x"02987058",
  1192 => x"486b87cc",
  1193 => x"a6c49872",
  1194 => x"05987058",
  1195 => x"7bc587f4",
  1196 => x"c148d4ff",
  1197 => x"78c378d3",
  1198 => x"9872486b",
  1199 => x"7058a6c4",
  1200 => x"87cc0298",
  1201 => x"9872486b",
  1202 => x"7058a6c4",
  1203 => x"87f40598",
  1204 => x"486b7bc4",
  1205 => x"a6c49872",
  1206 => x"02987058",
  1207 => x"486b87cc",
  1208 => x"a6c49872",
  1209 => x"05987058",
  1210 => x"d1c487f4",
  1211 => x"029d757b",
  1212 => x"c887f2c0",
  1213 => x"04adb7c0",
  1214 => x"8d4a87c4",
  1215 => x"4a7587c4",
  1216 => x"49724dc0",
  1217 => x"99718ac1",
  1218 => x"ff87ce02",
  1219 => x"78c048d4",
  1220 => x"8ac14972",
  1221 => x"f2059971",
  1222 => x"48d4ff87",
  1223 => x"757878c0",
  1224 => x"ceff059d",
  1225 => x"c0c0c887",
  1226 => x"72486b4a",
  1227 => x"58a6c498",
  1228 => x"cc029870",
  1229 => x"72486b87",
  1230 => x"58a6c498",
  1231 => x"f4059870",
  1232 => x"6b7bd087",
  1233 => x"c4987248",
  1234 => x"987058a6",
  1235 => x"6b87cc02",
  1236 => x"c4987248",
  1237 => x"987058a6",
  1238 => x"c587f405",
  1239 => x"48d4ff7b",
  1240 => x"c078d3c1",
  1241 => x"72486b78",
  1242 => x"58a6c498",
  1243 => x"cc029870",
  1244 => x"72486b87",
  1245 => x"58a6c498",
  1246 => x"f4059870",
  1247 => x"267bc487",
  1248 => x"0e87ecf6",
  1249 => x"5d5c5b5e",
  1250 => x"7186f40e",
  1251 => x"4cd0ff4d",
  1252 => x"4bc0c0c8",
  1253 => x"c0c31e75",
  1254 => x"e8e549d0",
  1255 => x"7086c487",
  1256 => x"c4c60298",
  1257 => x"d4c0c387",
  1258 => x"49757ebf",
  1259 => x"c887f7f6",
  1260 => x"1e7058a6",
  1261 => x"1e49a5c8",
  1262 => x"1ec0d5c1",
  1263 => x"87fcf2fe",
  1264 => x"486c86cc",
  1265 => x"a6cc9873",
  1266 => x"02987058",
  1267 => x"486c87cc",
  1268 => x"a6cc9873",
  1269 => x"05987058",
  1270 => x"7cc587f4",
  1271 => x"c148d4ff",
  1272 => x"c0c378d5",
  1273 => x"c149bfcc",
  1274 => x"4a66c481",
  1275 => x"32c68ac1",
  1276 => x"b0714872",
  1277 => x"7808d4ff",
  1278 => x"9873486c",
  1279 => x"7058a6cc",
  1280 => x"87cc0298",
  1281 => x"9873486c",
  1282 => x"7058a6c8",
  1283 => x"87f40598",
  1284 => x"d4ff7cc4",
  1285 => x"78ffc348",
  1286 => x"9873486c",
  1287 => x"7058a6c8",
  1288 => x"87cc0298",
  1289 => x"9873486c",
  1290 => x"7058a6c8",
  1291 => x"87f40598",
  1292 => x"d4ff7cc5",
  1293 => x"78d3c148",
  1294 => x"486c78c1",
  1295 => x"a6c89873",
  1296 => x"02987058",
  1297 => x"486c87cc",
  1298 => x"a6c89873",
  1299 => x"05987058",
  1300 => x"7cc487f4",
  1301 => x"d0c2026e",
  1302 => x"f4f2c287",
  1303 => x"c0c31e4d",
  1304 => x"c8e749d0",
  1305 => x"7086c487",
  1306 => x"87c50598",
  1307 => x"cac348c0",
  1308 => x"c8486e87",
  1309 => x"04a8b7c0",
  1310 => x"6e4a87cb",
  1311 => x"88c0c848",
  1312 => x"c458a6c4",
  1313 => x"c04a6e87",
  1314 => x"73486c7e",
  1315 => x"58a6c898",
  1316 => x"cc029870",
  1317 => x"73486c87",
  1318 => x"58a6c898",
  1319 => x"f4059870",
  1320 => x"ff7ccd87",
  1321 => x"d4c148d4",
  1322 => x"c1497278",
  1323 => x"0299718a",
  1324 => x"481587d0",
  1325 => x"7808d4ff",
  1326 => x"8ac14972",
  1327 => x"ff059971",
  1328 => x"486c87f0",
  1329 => x"a6c89873",
  1330 => x"02987058",
  1331 => x"486c87cd",
  1332 => x"a6c89873",
  1333 => x"05987058",
  1334 => x"c487f3ff",
  1335 => x"d0c0c37c",
  1336 => x"87e6e449",
  1337 => x"f0fd056e",
  1338 => x"73486c87",
  1339 => x"58a6c498",
  1340 => x"cd029870",
  1341 => x"73486c87",
  1342 => x"58a6c498",
  1343 => x"ff059870",
  1344 => x"7cc587f3",
  1345 => x"c148d4ff",
  1346 => x"78c078d3",
  1347 => x"9873486c",
  1348 => x"7058a6c4",
  1349 => x"87cd0298",
  1350 => x"9873486c",
  1351 => x"7058a6c4",
  1352 => x"f3ff0598",
  1353 => x"d07cc487",
  1354 => x"c11e7587",
  1355 => x"fe1ee6d5",
  1356 => x"c887c9ed",
  1357 => x"c248c086",
  1358 => x"f448c187",
  1359 => x"87efef8e",
  1360 => x"6e65704f",
  1361 => x"66206465",
  1362 => x"2c656c69",
  1363 => x"616f6c20",
  1364 => x"676e6964",
  1365 => x"2c732520",
  1366 => x"64692820",
  1367 => x"64252078",
  1368 => x"2e2e2e29",
  1369 => x"6143000a",
  1370 => x"2074276e",
  1371 => x"6e65706f",
  1372 => x"0a732520",
  1373 => x"6f6f4c00",
  1374 => x"676e696b",
  1375 => x"726f6620",
  1376 => x"6c696620",
  1377 => x"64252065",
  1378 => x"6946000a",
  1379 => x"2520656c",
  1380 => x"53000a73",
  1381 => x"63656c65",
  1382 => x"20646574",
  1383 => x"6d6f7266",
  1384 => x"20642520",
  1385 => x"6425202b",
  1386 => x"696c000a",
  1387 => x"6f727473",
  1388 => x"6b73206d",
  1389 => x"69707069",
  1390 => x"2520676e",
  1391 => x"64202c64",
  1392 => x"6e657269",
  1393 => x"65697274",
  1394 => x"64252073",
  1395 => x"80000a20",
  1396 => x"63614220",
  1397 => x"7573006b",
  1398 => x"6e656d62",
  1399 => x"61632075",
  1400 => x"61626c6c",
  1401 => x"4c006b63",
  1402 => x"2064616f",
  1403 => x"00202e2a",
  1404 => x"64616f4c",
  1405 => x"00203a00",
  1406 => x"6f636544",
  1407 => x"20646564",
  1408 => x"6f206425",
  1409 => x"6f697470",
  1410 => x"000a736e",
  1411 => x"65676150",
  1412 => x"0a642520",
  1413 => x"42208000",
  1414 => x"006b6361",
  1415 => x"78452080",
  1416 => x"4e007469",
  1417 => x"20747865",
  1418 => x"72616863",
  1419 => x"0a632520",
  1420 => x"78614d00",
  1421 => x"65676170",
  1422 => x"0a642520",
  1423 => x"4d4f5200",
  1424 => x"616f6c20",
  1425 => x"0a646564",
  1426 => x"4d4f5200",
  1427 => x"616f6c20",
  1428 => x"61662064",
  1429 => x"64656c69",
  1430 => x"6e49000a",
  1431 => x"61697469",
  1432 => x"697a696c",
  1433 => x"5320676e",
  1434 => x"61632044",
  1435 => x"000a6472",
  1436 => x"65766148",
  1437 => x"0a445320",
  1438 => x"5b5e0e00",
  1439 => x"1e0e5d5c",
  1440 => x"4cc04b71",
  1441 => x"d5c11e73",
  1442 => x"e7fe1ef5",
  1443 => x"86c887ee",
  1444 => x"abb74dc0",
  1445 => x"87e9c004",
  1446 => x"1ee6c5c1",
  1447 => x"c4029d75",
  1448 => x"c24ac087",
  1449 => x"724ac187",
  1450 => x"87fee049",
  1451 => x"58a686c4",
  1452 => x"056e84c1",
  1453 => x"4c7387c2",
  1454 => x"b77385c1",
  1455 => x"d7ff06ac",
  1456 => x"26486e87",
  1457 => x"0e87e8e9",
  1458 => x"5d5c5b5e",
  1459 => x"1e4c710e",
  1460 => x"bfdcc0c3",
  1461 => x"d3d6c11e",
  1462 => x"dfe6fe1e",
  1463 => x"dcc0c387",
  1464 => x"817449bf",
  1465 => x"7087d2fe",
  1466 => x"d6c11e4d",
  1467 => x"e6fe1eca",
  1468 => x"86d487ca",
  1469 => x"d3029d75",
  1470 => x"c4fbc287",
  1471 => x"cb4a754b",
  1472 => x"c6ebfe49",
  1473 => x"c4fbc287",
  1474 => x"87f7f149",
  1475 => x"49fdfbc1",
  1476 => x"87c6c7c1",
  1477 => x"87e2c7c1",
  1478 => x"1e87d4e8",
  1479 => x"4b711e73",
  1480 => x"dcc0c349",
  1481 => x"d0fd81bf",
  1482 => x"9a4a7087",
  1483 => x"4987c502",
  1484 => x"87f3dcff",
  1485 => x"48dcc0c3",
  1486 => x"497378c0",
  1487 => x"e787e9c1",
  1488 => x"731e87f1",
  1489 => x"c44b711e",
  1490 => x"c1024aa3",
  1491 => x"8ac187c8",
  1492 => x"8a87dc02",
  1493 => x"87f1c002",
  1494 => x"c4c1058a",
  1495 => x"dcc0c387",
  1496 => x"fcc002bf",
  1497 => x"88c14887",
  1498 => x"58e0c0c3",
  1499 => x"c387f2c0",
  1500 => x"49bfdcc0",
  1501 => x"c0c389d0",
  1502 => x"b7c059e0",
  1503 => x"e0c003a9",
  1504 => x"dcc0c387",
  1505 => x"d878c048",
  1506 => x"dcc0c387",
  1507 => x"80c148bf",
  1508 => x"58e0c0c3",
  1509 => x"c0c387cb",
  1510 => x"d048bfdc",
  1511 => x"e0c0c380",
  1512 => x"c3497358",
  1513 => x"87cbe687",
  1514 => x"5c5b5e0e",
  1515 => x"86f00e5d",
  1516 => x"c259a6d0",
  1517 => x"c04df4f2",
  1518 => x"c0fbc24c",
  1519 => x"c0c31ebf",
  1520 => x"c11ebfdc",
  1521 => x"fe1eead6",
  1522 => x"cc87f1e2",
  1523 => x"48a6c486",
  1524 => x"c0c378c0",
  1525 => x"c048bfdc",
  1526 => x"c106a8b7",
  1527 => x"f2c287c2",
  1528 => x"029848f4",
  1529 => x"c187f9c0",
  1530 => x"c81ee6c5",
  1531 => x"87c70266",
  1532 => x"c048a6c4",
  1533 => x"c487c578",
  1534 => x"78c148a6",
  1535 => x"ff4966c4",
  1536 => x"c487e7db",
  1537 => x"c14d7086",
  1538 => x"4866c484",
  1539 => x"a6c880c1",
  1540 => x"dcc0c358",
  1541 => x"03acb7bf",
  1542 => x"9d7587c6",
  1543 => x"87c7ff05",
  1544 => x"9d754cc0",
  1545 => x"87e5c302",
  1546 => x"1ee6c5c1",
  1547 => x"c70266c8",
  1548 => x"48a6cc87",
  1549 => x"87c578c0",
  1550 => x"c148a6cc",
  1551 => x"4966cc78",
  1552 => x"87e6daff",
  1553 => x"58a686c4",
  1554 => x"ecc2026e",
  1555 => x"81cb4987",
  1556 => x"d0496997",
  1557 => x"d9c10299",
  1558 => x"dbdcc187",
  1559 => x"cc49744b",
  1560 => x"fdfbc191",
  1561 => x"4aa1c881",
  1562 => x"81c17a73",
  1563 => x"7451ffc3",
  1564 => x"c391de49",
  1565 => x"714df0c0",
  1566 => x"97c1c285",
  1567 => x"49a5c17d",
  1568 => x"c251e0c0",
  1569 => x"bf97c4fb",
  1570 => x"c187d202",
  1571 => x"4ba5c284",
  1572 => x"4ac4fbc2",
  1573 => x"e4fe49db",
  1574 => x"dcc187f1",
  1575 => x"49a5cd87",
  1576 => x"84c151c0",
  1577 => x"6e4ba5c2",
  1578 => x"fe49cb4a",
  1579 => x"c187dce4",
  1580 => x"497487c7",
  1581 => x"fbc191cc",
  1582 => x"81c881fd",
  1583 => x"79c7dbc1",
  1584 => x"97c4fbc2",
  1585 => x"87d902bf",
  1586 => x"91de4974",
  1587 => x"c0c384c1",
  1588 => x"83714bf0",
  1589 => x"4ac4fbc2",
  1590 => x"e3fe49dd",
  1591 => x"d8c087ed",
  1592 => x"de4b7487",
  1593 => x"f0c0c393",
  1594 => x"49a3cb83",
  1595 => x"84c151c0",
  1596 => x"cb4a6e73",
  1597 => x"d2e3fe49",
  1598 => x"4866c487",
  1599 => x"a6c880c1",
  1600 => x"acb7c758",
  1601 => x"87c5c003",
  1602 => x"dbfc056e",
  1603 => x"acb7c787",
  1604 => x"87d3c003",
  1605 => x"91de4974",
  1606 => x"81f0c0c3",
  1607 => x"84c151c0",
  1608 => x"04acb7c7",
  1609 => x"c187edff",
  1610 => x"c048d2fd",
  1611 => x"d1fdc150",
  1612 => x"c150c248",
  1613 => x"c148d9fd",
  1614 => x"c178e6e5",
  1615 => x"c148d5fd",
  1616 => x"c178cfd7",
  1617 => x"c148e5fd",
  1618 => x"cc78c2dd",
  1619 => x"fac04966",
  1620 => x"8ef087c9",
  1621 => x"87d7dfff",
  1622 => x"c34a711e",
  1623 => x"725ad0c0",
  1624 => x"87c4f949",
  1625 => x"731e4f26",
  1626 => x"494b711e",
  1627 => x"fbc191cc",
  1628 => x"81c181fd",
  1629 => x"c0c34811",
  1630 => x"d7c158cc",
  1631 => x"e0fe49d6",
  1632 => x"f0c087e5",
  1633 => x"e1fe49a3",
  1634 => x"49c087d1",
  1635 => x"ff87f8d2",
  1636 => x"0e87e0de",
  1637 => x"5d5c5b5e",
  1638 => x"7186f00e",
  1639 => x"91cc494c",
  1640 => x"81fdfbc1",
  1641 => x"c47ea1c3",
  1642 => x"c0c348a6",
  1643 => x"6e78bfc4",
  1644 => x"c44abf97",
  1645 => x"2b724b66",
  1646 => x"124aa1c1",
  1647 => x"58a6cc48",
  1648 => x"83c19b70",
  1649 => x"699781c2",
  1650 => x"04abb749",
  1651 => x"4bc087c2",
  1652 => x"4abf976e",
  1653 => x"724966c8",
  1654 => x"c4b9ff31",
  1655 => x"4d739966",
  1656 => x"b5713572",
  1657 => x"5dc8c0c3",
  1658 => x"c348d4ff",
  1659 => x"d0ff78ff",
  1660 => x"c0c848bf",
  1661 => x"a6d098c0",
  1662 => x"02987058",
  1663 => x"d0ff87d0",
  1664 => x"c0c848bf",
  1665 => x"a6c498c0",
  1666 => x"05987058",
  1667 => x"d0ff87f0",
  1668 => x"78e1c048",
  1669 => x"de48d4ff",
  1670 => x"7d0d7078",
  1671 => x"c848750d",
  1672 => x"d4ff28b7",
  1673 => x"48757808",
  1674 => x"ff28b7d0",
  1675 => x"757808d4",
  1676 => x"28b7d848",
  1677 => x"7808d4ff",
  1678 => x"48bfd0ff",
  1679 => x"98c0c0c8",
  1680 => x"7058a6c4",
  1681 => x"87d00298",
  1682 => x"48bfd0ff",
  1683 => x"98c0c0c8",
  1684 => x"7058a6c4",
  1685 => x"87f00598",
  1686 => x"c048d0ff",
  1687 => x"1ec778e0",
  1688 => x"fbc11ec0",
  1689 => x"c0c31efd",
  1690 => x"cc49bfc8",
  1691 => x"c0497487",
  1692 => x"e487e8f5",
  1693 => x"f6daff8e",
  1694 => x"5b5e0e87",
  1695 => x"ff0e5d5c",
  1696 => x"a6d886d8",
  1697 => x"48a6c859",
  1698 => x"80c478c0",
  1699 => x"80c478c0",
  1700 => x"d4ff78c0",
  1701 => x"78ffc348",
  1702 => x"48bfd0ff",
  1703 => x"98c0c0c8",
  1704 => x"7058a6c4",
  1705 => x"87d00298",
  1706 => x"48bfd0ff",
  1707 => x"98c0c0c8",
  1708 => x"7058a6c4",
  1709 => x"87f00598",
  1710 => x"c048d0ff",
  1711 => x"d4ff78e1",
  1712 => x"ff78d448",
  1713 => x"ff87dfd7",
  1714 => x"ffc348d4",
  1715 => x"1e4d6878",
  1716 => x"1ee3d8c1",
  1717 => x"87e4d6fe",
  1718 => x"fbc086c8",
  1719 => x"c5c102ad",
  1720 => x"66f8c087",
  1721 => x"6a82c44a",
  1722 => x"c11e727e",
  1723 => x"c448e7d7",
  1724 => x"a1c84966",
  1725 => x"7141204a",
  1726 => x"87f905aa",
  1727 => x"4a265110",
  1728 => x"4966f8c0",
  1729 => x"e5c181c8",
  1730 => x"496a79d8",
  1731 => x"0d7181c8",
  1732 => x"c10d7d97",
  1733 => x"6a1ed81e",
  1734 => x"ff81c849",
  1735 => x"c887ded6",
  1736 => x"48a6d086",
  1737 => x"9d7578c1",
  1738 => x"87e8c902",
  1739 => x"c14866d0",
  1740 => x"a8b766c0",
  1741 => x"87dcc903",
  1742 => x"c348d4ff",
  1743 => x"486878ff",
  1744 => x"c488c6c1",
  1745 => x"987058a6",
  1746 => x"4887db02",
  1747 => x"a6c488c9",
  1748 => x"02987058",
  1749 => x"4887ebc3",
  1750 => x"a6c488c1",
  1751 => x"02987058",
  1752 => x"c887c5c1",
  1753 => x"66d487d6",
  1754 => x"87f3c005",
  1755 => x"cc4966d0",
  1756 => x"66f8c091",
  1757 => x"4aa1c481",
  1758 => x"1e717e6a",
  1759 => x"48f0d7c1",
  1760 => x"c44966c4",
  1761 => x"41204aa1",
  1762 => x"f905aa71",
  1763 => x"26511087",
  1764 => x"c181c849",
  1765 => x"d079d8e5",
  1766 => x"80c14866",
  1767 => x"ff58a6d4",
  1768 => x"7087c3d4",
  1769 => x"87dac74d",
  1770 => x"87cbd6ff",
  1771 => x"7058a6cc",
  1772 => x"ccd8c11e",
  1773 => x"c3d3fe1e",
  1774 => x"6686c887",
  1775 => x"b766cc48",
  1776 => x"87c606a8",
  1777 => x"c848a6cc",
  1778 => x"d5ff7866",
  1779 => x"ecc087e9",
  1780 => x"edc105a8",
  1781 => x"0566d487",
  1782 => x"d087dec1",
  1783 => x"91cc4966",
  1784 => x"8166f8c0",
  1785 => x"6a4aa1c4",
  1786 => x"4aa1c14c",
  1787 => x"c25266c8",
  1788 => x"81c87997",
  1789 => x"79e6e5c1",
  1790 => x"c348d4ff",
  1791 => x"4d6878ff",
  1792 => x"e0c0029d",
  1793 => x"adfbc087",
  1794 => x"7487da02",
  1795 => x"0d7d970d",
  1796 => x"d4ff84c1",
  1797 => x"78ffc348",
  1798 => x"029d4d68",
  1799 => x"fbc087c7",
  1800 => x"e6ff05ad",
  1801 => x"54e0c087",
  1802 => x"c054c1c2",
  1803 => x"66d07c97",
  1804 => x"d480c148",
  1805 => x"c9c558a6",
  1806 => x"e9d1ff87",
  1807 => x"c54d7087",
  1808 => x"66c887c0",
  1809 => x"a866d448",
  1810 => x"87e7c405",
  1811 => x"c048a6d8",
  1812 => x"e2d3ff78",
  1813 => x"a6e0c087",
  1814 => x"dad3ff58",
  1815 => x"a6e4c087",
  1816 => x"a8ecc058",
  1817 => x"87cac005",
  1818 => x"48a6e0c0",
  1819 => x"c07866dc",
  1820 => x"d4ff87c6",
  1821 => x"78ffc348",
  1822 => x"cc4966d0",
  1823 => x"66f8c091",
  1824 => x"c4807148",
  1825 => x"496e58a6",
  1826 => x"66dc81c3",
  1827 => x"66e0c051",
  1828 => x"dc81c149",
  1829 => x"48c18966",
  1830 => x"49703071",
  1831 => x"4a6e89c1",
  1832 => x"097282c1",
  1833 => x"6e097997",
  1834 => x"6e50c248",
  1835 => x"c181c849",
  1836 => x"c379d3e6",
  1837 => x"49bfc4c0",
  1838 => x"29b766dc",
  1839 => x"484a6a97",
  1840 => x"e8c09871",
  1841 => x"486e58a6",
  1842 => x"a6c880c4",
  1843 => x"bf66c458",
  1844 => x"4866d44c",
  1845 => x"02a866c8",
  1846 => x"dc87c8c0",
  1847 => x"78c048a6",
  1848 => x"dc87c5c0",
  1849 => x"78c148a6",
  1850 => x"c01e66dc",
  1851 => x"49741ee0",
  1852 => x"87c9cfff",
  1853 => x"4d7086c8",
  1854 => x"06adb7c0",
  1855 => x"7587d5c1",
  1856 => x"bf66c484",
  1857 => x"81e0c049",
  1858 => x"c14b8974",
  1859 => x"714af5d7",
  1860 => x"87f7d2fe",
  1861 => x"66d884c2",
  1862 => x"dc80c148",
  1863 => x"e4c058a6",
  1864 => x"81c14966",
  1865 => x"c002a970",
  1866 => x"a6dc87c8",
  1867 => x"c078c048",
  1868 => x"a6dc87c5",
  1869 => x"dc78c148",
  1870 => x"66c81e66",
  1871 => x"e0c049bf",
  1872 => x"71897481",
  1873 => x"ff49741e",
  1874 => x"c887f2cd",
  1875 => x"a8b7c086",
  1876 => x"87c2ff01",
  1877 => x"c11e66d8",
  1878 => x"fe1ef8d7",
  1879 => x"c887ddcc",
  1880 => x"c2496e86",
  1881 => x"5166d881",
  1882 => x"c14866d0",
  1883 => x"58a6d480",
  1884 => x"ff87cfc0",
  1885 => x"7087efcc",
  1886 => x"87c6c04d",
  1887 => x"87e6ccff",
  1888 => x"9d754d70",
  1889 => x"87ccc002",
  1890 => x"c14866d0",
  1891 => x"a8b766c0",
  1892 => x"87e4f604",
  1893 => x"c74866d0",
  1894 => x"c003a8b7",
  1895 => x"66d087e3",
  1896 => x"c091cc49",
  1897 => x"c48166f8",
  1898 => x"4a6a4aa1",
  1899 => x"81c852c0",
  1900 => x"66d079c0",
  1901 => x"d480c148",
  1902 => x"b7c758a6",
  1903 => x"ddff04a8",
  1904 => x"0266d487",
  1905 => x"c087ebc0",
  1906 => x"c14966f8",
  1907 => x"f8c081d4",
  1908 => x"d5c14a66",
  1909 => x"c252c082",
  1910 => x"66f8c051",
  1911 => x"81dcc149",
  1912 => x"79e6e5c1",
  1913 => x"4966f8c0",
  1914 => x"c181d8c1",
  1915 => x"c079d5d8",
  1916 => x"f8c087d6",
  1917 => x"d8c14966",
  1918 => x"dcd8c181",
  1919 => x"66f8c079",
  1920 => x"81dcc149",
  1921 => x"79fae3c2",
  1922 => x"c11e66cc",
  1923 => x"fe1ef1d8",
  1924 => x"c887e9c9",
  1925 => x"bfd0ff86",
  1926 => x"c0c0c848",
  1927 => x"58a6c498",
  1928 => x"c0029870",
  1929 => x"d0ff87d1",
  1930 => x"c0c848bf",
  1931 => x"a6c498c0",
  1932 => x"05987058",
  1933 => x"ff87efff",
  1934 => x"e0c048d0",
  1935 => x"4866cc78",
  1936 => x"ff8ed8ff",
  1937 => x"1e87e8cb",
  1938 => x"1ec01ec7",
  1939 => x"1efdfbc1",
  1940 => x"bfc8c0c3",
  1941 => x"87e1f049",
  1942 => x"49fdfbc1",
  1943 => x"87fae9c0",
  1944 => x"4f268ef4",
  1945 => x"ca1e731e",
  1946 => x"c0c387f4",
  1947 => x"50c048e0",
  1948 => x"c348d4ff",
  1949 => x"d9c178ff",
  1950 => x"ccfe49da",
  1951 => x"d9fe87e9",
  1952 => x"987087e5",
  1953 => x"fe87cd02",
  1954 => x"7087e5e6",
  1955 => x"87c40298",
  1956 => x"87c24bc1",
  1957 => x"9b734bc0",
  1958 => x"c187c802",
  1959 => x"fe49f0d9",
  1960 => x"c387c4cc",
  1961 => x"c048c8c0",
  1962 => x"dafe4978",
  1963 => x"87dac487",
  1964 => x"c087ffc9",
  1965 => x"c587fdec",
  1966 => x"87c0ce49",
  1967 => x"c4029870",
  1968 => x"feceff87",
  1969 => x"49f8c187",
  1970 => x"7087f1cd",
  1971 => x"dfff0298",
  1972 => x"029b7387",
  1973 => x"c0c387d8",
  1974 => x"d2ff49e0",
  1975 => x"987087e5",
  1976 => x"c187cb02",
  1977 => x"fe49fdd8",
  1978 => x"ff87fcca",
  1979 => x"d9c187c2",
  1980 => x"cafe49c9",
  1981 => x"f7fe87f1",
  1982 => x"f6c8ff87",
  1983 => x"00000287",
  1984 => x"00303000",
  1985 => x"0016c700",
  1986 => x"00000200",
  1987 => x"00304e00",
  1988 => x"0016c700",
  1989 => x"00000200",
  1990 => x"00306c00",
  1991 => x"0016c700",
  1992 => x"00000200",
  1993 => x"00308a00",
  1994 => x"0016c700",
  1995 => x"00000200",
  1996 => x"0030a800",
  1997 => x"0016c700",
  1998 => x"00000200",
  1999 => x"0030c600",
  2000 => x"0016c700",
  2001 => x"00000200",
  2002 => x"0030e400",
  2003 => x"0016c700",
  2004 => x"00000200",
  2005 => x"00000000",
  2006 => x"00196600",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00174200",
  2010 => x"c11e1e00",
  2011 => x"a6c487d5",
  2012 => x"4f262658",
  2013 => x"fe4a711e",
  2014 => x"78c048f0",
  2015 => x"0a7a0acd",
  2016 => x"49cafec1",
  2017 => x"87dfc8fe",
  2018 => x"65534f26",
  2019 => x"61682074",
  2020 => x"656c646e",
  2021 => x"49000a72",
  2022 => x"6e69206e",
  2023 => x"72726574",
  2024 => x"20747075",
  2025 => x"736e6f63",
  2026 => x"63757274",
  2027 => x"0a726f74",
  2028 => x"fec11e00",
  2029 => x"c7fe49d7",
  2030 => x"fdc187ed",
  2031 => x"f3fe49e9",
  2032 => x"1e4f2687",
  2033 => x"48bff0fe",
  2034 => x"fe1e4f26",
  2035 => x"78c148f0",
  2036 => x"fe1e4f26",
  2037 => x"78c048f0",
  2038 => x"711e4f26",
  2039 => x"c47ac04a",
  2040 => x"79c049a2",
  2041 => x"c049a2c8",
  2042 => x"49a2cc79",
  2043 => x"4f2679c0",
  2044 => x"5c5b5e0e",
  2045 => x"7186f80e",
  2046 => x"49a4c84c",
  2047 => x"6b4ba4cc",
  2048 => x"c480c148",
  2049 => x"98cf58a6",
  2050 => x"6958a6c8",
  2051 => x"a866c448",
  2052 => x"6b87d405",
  2053 => x"c480c148",
  2054 => x"98cf58a6",
  2055 => x"6958a6c8",
  2056 => x"a866c448",
  2057 => x"fe87ec02",
  2058 => x"d0c187e8",
  2059 => x"486b49a4",
  2060 => x"a6c490c4",
  2061 => x"d4817058",
  2062 => x"486b7966",
  2063 => x"a6c880c1",
  2064 => x"7098cf58",
  2065 => x"87d2c17b",
  2066 => x"f887fffd",
  2067 => x"2687c28e",
  2068 => x"264c264d",
  2069 => x"0e4f264b",
  2070 => x"5d5c5b5e",
  2071 => x"7186f80e",
  2072 => x"4ca5c44d",
  2073 => x"a86c486d",
  2074 => x"ff87c505",
  2075 => x"87e5c048",
  2076 => x"d087dffd",
  2077 => x"486c4ba5",
  2078 => x"a6c490c4",
  2079 => x"6b837058",
  2080 => x"9bffc34b",
  2081 => x"80c1486c",
  2082 => x"cf58a6c8",
  2083 => x"fc7c7098",
  2084 => x"497387f8",
  2085 => x"fe8ef848",
  2086 => x"731e87f5",
  2087 => x"fc86f81e",
  2088 => x"bfe087f0",
  2089 => x"e0c0494b",
  2090 => x"c00299c0",
  2091 => x"4a7387e7",
  2092 => x"c39affc3",
  2093 => x"48bfc2c4",
  2094 => x"a6c490c4",
  2095 => x"d2c4c358",
  2096 => x"72817049",
  2097 => x"c2c4c379",
  2098 => x"80c148bf",
  2099 => x"cf58a6c8",
  2100 => x"c6c4c398",
  2101 => x"d0497358",
  2102 => x"c00299c0",
  2103 => x"c4c387f2",
  2104 => x"c348bfca",
  2105 => x"a8bfcec4",
  2106 => x"87e4c002",
  2107 => x"bfcac4c3",
  2108 => x"c490c448",
  2109 => x"c5c358a6",
  2110 => x"817049d2",
  2111 => x"786948e0",
  2112 => x"bfcac4c3",
  2113 => x"c880c148",
  2114 => x"98cf58a6",
  2115 => x"58cec4c3",
  2116 => x"c487f0fa",
  2117 => x"f1fa58a6",
  2118 => x"fc8ef887",
  2119 => x"c31e87f5",
  2120 => x"fa49c2c4",
  2121 => x"c2c287f4",
  2122 => x"c7f949da",
  2123 => x"87f5c387",
  2124 => x"731e4f26",
  2125 => x"c2c4c31e",
  2126 => x"87dbfc49",
  2127 => x"b7c04a70",
  2128 => x"ccc204aa",
  2129 => x"aaf0c387",
  2130 => x"c287c905",
  2131 => x"c148ddc7",
  2132 => x"87edc178",
  2133 => x"05aae0c3",
  2134 => x"c7c287c9",
  2135 => x"78c148e1",
  2136 => x"c287dec1",
  2137 => x"02bfe1c7",
  2138 => x"c0c287c6",
  2139 => x"87c24ba2",
  2140 => x"c7c24b72",
  2141 => x"c002bfdd",
  2142 => x"497387e0",
  2143 => x"9129b7c4",
  2144 => x"81e5c7c2",
  2145 => x"9acf4a73",
  2146 => x"48c192c2",
  2147 => x"4a703072",
  2148 => x"4872baff",
  2149 => x"79709869",
  2150 => x"497387db",
  2151 => x"9129b7c4",
  2152 => x"81e5c7c2",
  2153 => x"9acf4a73",
  2154 => x"48c392c2",
  2155 => x"4a703072",
  2156 => x"70b06948",
  2157 => x"e1c7c279",
  2158 => x"c278c048",
  2159 => x"c048ddc7",
  2160 => x"c2c4c378",
  2161 => x"87cffa49",
  2162 => x"b7c04a70",
  2163 => x"f4fd03aa",
  2164 => x"c448c087",
  2165 => x"264d2687",
  2166 => x"264b264c",
  2167 => x"0000004f",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"4ac01e00",
  2186 => x"91c44972",
  2187 => x"81e5c7c2",
  2188 => x"82c179c0",
  2189 => x"04aab7d0",
  2190 => x"4f2687ee",
  2191 => x"5c5b5e0e",
  2192 => x"4d710e5d",
  2193 => x"7587cbf6",
  2194 => x"2ab7c44a",
  2195 => x"e5c7c292",
  2196 => x"cf4c7582",
  2197 => x"6a94c29c",
  2198 => x"2b744b49",
  2199 => x"48c29bc3",
  2200 => x"4c703074",
  2201 => x"4874bcff",
  2202 => x"7a709871",
  2203 => x"7387dbf5",
  2204 => x"87e1fd48",
  2205 => x"d0ff1e1e",
  2206 => x"c0c848bf",
  2207 => x"a6c498c0",
  2208 => x"02987058",
  2209 => x"d0ff87d0",
  2210 => x"c0c848bf",
  2211 => x"a6c498c0",
  2212 => x"05987058",
  2213 => x"d0ff87f0",
  2214 => x"78e1c448",
  2215 => x"d4ff4871",
  2216 => x"66c87808",
  2217 => x"08d4ff48",
  2218 => x"4f262678",
  2219 => x"4a711e1e",
  2220 => x"1e4966c8",
  2221 => x"fbfe4972",
  2222 => x"ff86c487",
  2223 => x"c848bfd0",
  2224 => x"c498c0c0",
  2225 => x"987058a6",
  2226 => x"ff87d002",
  2227 => x"c848bfd0",
  2228 => x"c498c0c0",
  2229 => x"987058a6",
  2230 => x"ff87f005",
  2231 => x"e0c048d0",
  2232 => x"4f262678",
  2233 => x"711e731e",
  2234 => x"1e66c84b",
  2235 => x"e0c14a73",
  2236 => x"f7fe49a2",
  2237 => x"87c42687",
  2238 => x"4c264d26",
  2239 => x"4f264b26",
  2240 => x"d0ff1e1e",
  2241 => x"c0c848bf",
  2242 => x"a6c498c0",
  2243 => x"02987058",
  2244 => x"d0ff87d0",
  2245 => x"c0c848bf",
  2246 => x"a6c498c0",
  2247 => x"05987058",
  2248 => x"d0ff87f0",
  2249 => x"78c9c448",
  2250 => x"d4ff4871",
  2251 => x"26267808",
  2252 => x"711e1e4f",
  2253 => x"c7ff494a",
  2254 => x"bfd0ff87",
  2255 => x"c0c0c848",
  2256 => x"58a6c498",
  2257 => x"d0029870",
  2258 => x"bfd0ff87",
  2259 => x"c0c0c848",
  2260 => x"58a6c498",
  2261 => x"f0059870",
  2262 => x"48d0ff87",
  2263 => x"262678c8",
  2264 => x"1e731e4f",
  2265 => x"c34b711e",
  2266 => x"02bfdec6",
  2267 => x"ccc387c3",
  2268 => x"bfd0ff87",
  2269 => x"c0c0c848",
  2270 => x"58a6c498",
  2271 => x"d0029870",
  2272 => x"bfd0ff87",
  2273 => x"c0c0c848",
  2274 => x"58a6c498",
  2275 => x"f0059870",
  2276 => x"48d0ff87",
  2277 => x"7378c9c4",
  2278 => x"b0e0c048",
  2279 => x"7808d4ff",
  2280 => x"48d2c6c3",
  2281 => x"66cc78c0",
  2282 => x"c387c502",
  2283 => x"87c249ff",
  2284 => x"c6c349c0",
  2285 => x"66d059da",
  2286 => x"c587c602",
  2287 => x"c44ad5d5",
  2288 => x"ffffcf87",
  2289 => x"dec6c34a",
  2290 => x"dec6c35a",
  2291 => x"2678c148",
  2292 => x"4d2687c4",
  2293 => x"4b264c26",
  2294 => x"5e0e4f26",
  2295 => x"0e5d5c5b",
  2296 => x"c6c34a71",
  2297 => x"724cbfda",
  2298 => x"87cb029a",
  2299 => x"c291c849",
  2300 => x"714bdbce",
  2301 => x"c287c483",
  2302 => x"c04bdbd2",
  2303 => x"7449134d",
  2304 => x"d6c6c399",
  2305 => x"b87148bf",
  2306 => x"7808d4ff",
  2307 => x"852cb7c1",
  2308 => x"04adb7c8",
  2309 => x"c6c387e7",
  2310 => x"c848bfd2",
  2311 => x"d6c6c380",
  2312 => x"87eefe58",
  2313 => x"711e731e",
  2314 => x"9a4a134b",
  2315 => x"7287cb02",
  2316 => x"87e6fe49",
  2317 => x"059a4a13",
  2318 => x"d9fe87f5",
  2319 => x"c31e1e87",
  2320 => x"49bfd2c6",
  2321 => x"48d2c6c3",
  2322 => x"c478a1c1",
  2323 => x"03a9b7c0",
  2324 => x"d4ff87db",
  2325 => x"d6c6c348",
  2326 => x"c6c378bf",
  2327 => x"c349bfd2",
  2328 => x"c148d2c6",
  2329 => x"c0c478a1",
  2330 => x"e504a9b7",
  2331 => x"bfd0ff87",
  2332 => x"c0c0c848",
  2333 => x"58a6c498",
  2334 => x"d0029870",
  2335 => x"bfd0ff87",
  2336 => x"c0c0c848",
  2337 => x"58a6c498",
  2338 => x"f0059870",
  2339 => x"48d0ff87",
  2340 => x"c6c378c8",
  2341 => x"78c048de",
  2342 => x"004f2626",
  2343 => x"00000000",
  2344 => x"00000000",
  2345 => x"5f5f0000",
  2346 => x"00000000",
  2347 => x"03000303",
  2348 => x"14000003",
  2349 => x"7f147f7f",
  2350 => x"0000147f",
  2351 => x"6b6b2e24",
  2352 => x"4c00123a",
  2353 => x"6c18366a",
  2354 => x"30003256",
  2355 => x"77594f7e",
  2356 => x"0040683a",
  2357 => x"03070400",
  2358 => x"00000000",
  2359 => x"633e1c00",
  2360 => x"00000041",
  2361 => x"3e634100",
  2362 => x"0800001c",
  2363 => x"1c1c3e2a",
  2364 => x"00082a3e",
  2365 => x"3e3e0808",
  2366 => x"00000808",
  2367 => x"60e08000",
  2368 => x"00000000",
  2369 => x"08080808",
  2370 => x"00000808",
  2371 => x"60600000",
  2372 => x"40000000",
  2373 => x"0c183060",
  2374 => x"00010306",
  2375 => x"4d597f3e",
  2376 => x"00003e7f",
  2377 => x"7f7f0604",
  2378 => x"00000000",
  2379 => x"59716342",
  2380 => x"0000464f",
  2381 => x"49496322",
  2382 => x"1800367f",
  2383 => x"7f13161c",
  2384 => x"0000107f",
  2385 => x"45456727",
  2386 => x"0000397d",
  2387 => x"494b7e3c",
  2388 => x"00003079",
  2389 => x"79710101",
  2390 => x"0000070f",
  2391 => x"49497f36",
  2392 => x"0000367f",
  2393 => x"69494f06",
  2394 => x"00001e3f",
  2395 => x"66660000",
  2396 => x"00000000",
  2397 => x"66e68000",
  2398 => x"00000000",
  2399 => x"14140808",
  2400 => x"00002222",
  2401 => x"14141414",
  2402 => x"00001414",
  2403 => x"14142222",
  2404 => x"00000808",
  2405 => x"59510302",
  2406 => x"3e00060f",
  2407 => x"555d417f",
  2408 => x"00001e1f",
  2409 => x"09097f7e",
  2410 => x"00007e7f",
  2411 => x"49497f7f",
  2412 => x"0000367f",
  2413 => x"41633e1c",
  2414 => x"00004141",
  2415 => x"63417f7f",
  2416 => x"00001c3e",
  2417 => x"49497f7f",
  2418 => x"00004141",
  2419 => x"09097f7f",
  2420 => x"00000101",
  2421 => x"49417f3e",
  2422 => x"00007a7b",
  2423 => x"08087f7f",
  2424 => x"00007f7f",
  2425 => x"7f7f4100",
  2426 => x"00000041",
  2427 => x"40406020",
  2428 => x"7f003f7f",
  2429 => x"361c087f",
  2430 => x"00004163",
  2431 => x"40407f7f",
  2432 => x"7f004040",
  2433 => x"060c067f",
  2434 => x"7f007f7f",
  2435 => x"180c067f",
  2436 => x"00007f7f",
  2437 => x"41417f3e",
  2438 => x"00003e7f",
  2439 => x"09097f7f",
  2440 => x"3e00060f",
  2441 => x"7f61417f",
  2442 => x"0000407e",
  2443 => x"19097f7f",
  2444 => x"0000667f",
  2445 => x"594d6f26",
  2446 => x"0000327b",
  2447 => x"7f7f0101",
  2448 => x"00000101",
  2449 => x"40407f3f",
  2450 => x"00003f7f",
  2451 => x"70703f0f",
  2452 => x"7f000f3f",
  2453 => x"3018307f",
  2454 => x"41007f7f",
  2455 => x"1c1c3663",
  2456 => x"01416336",
  2457 => x"7c7c0603",
  2458 => x"61010306",
  2459 => x"474d5971",
  2460 => x"00004143",
  2461 => x"417f7f00",
  2462 => x"01000041",
  2463 => x"180c0603",
  2464 => x"00406030",
  2465 => x"7f414100",
  2466 => x"0800007f",
  2467 => x"0603060c",
  2468 => x"8000080c",
  2469 => x"80808080",
  2470 => x"00008080",
  2471 => x"07030000",
  2472 => x"00000004",
  2473 => x"54547420",
  2474 => x"0000787c",
  2475 => x"44447f7f",
  2476 => x"0000387c",
  2477 => x"44447c38",
  2478 => x"00000044",
  2479 => x"44447c38",
  2480 => x"00007f7f",
  2481 => x"54547c38",
  2482 => x"0000185c",
  2483 => x"057f7e04",
  2484 => x"00000005",
  2485 => x"a4a4bc18",
  2486 => x"00007cfc",
  2487 => x"04047f7f",
  2488 => x"0000787c",
  2489 => x"7d3d0000",
  2490 => x"00000040",
  2491 => x"fd808080",
  2492 => x"0000007d",
  2493 => x"38107f7f",
  2494 => x"0000446c",
  2495 => x"7f3f0000",
  2496 => x"7c000040",
  2497 => x"0c180c7c",
  2498 => x"0000787c",
  2499 => x"04047c7c",
  2500 => x"0000787c",
  2501 => x"44447c38",
  2502 => x"0000387c",
  2503 => x"2424fcfc",
  2504 => x"0000183c",
  2505 => x"24243c18",
  2506 => x"0000fcfc",
  2507 => x"04047c7c",
  2508 => x"0000080c",
  2509 => x"54545c48",
  2510 => x"00002074",
  2511 => x"447f3f04",
  2512 => x"00000044",
  2513 => x"40407c3c",
  2514 => x"00007c7c",
  2515 => x"60603c1c",
  2516 => x"3c001c3c",
  2517 => x"6030607c",
  2518 => x"44003c7c",
  2519 => x"3810386c",
  2520 => x"0000446c",
  2521 => x"60e0bc1c",
  2522 => x"00001c3c",
  2523 => x"5c746444",
  2524 => x"0000444c",
  2525 => x"773e0808",
  2526 => x"00004141",
  2527 => x"7f7f0000",
  2528 => x"00000000",
  2529 => x"3e774141",
  2530 => x"02000808",
  2531 => x"02030101",
  2532 => x"7f000102",
  2533 => x"7f7f7f7f",
  2534 => x"08007f7f",
  2535 => x"3e1c1c08",
  2536 => x"7f7f7f3e",
  2537 => x"1c3e3e7f",
  2538 => x"0008081c",
  2539 => x"7c7c1810",
  2540 => x"00001018",
  2541 => x"7c7c3010",
  2542 => x"10001030",
  2543 => x"78606030",
  2544 => x"4200061e",
  2545 => x"3c183c66",
  2546 => x"78004266",
  2547 => x"c6c26a38",
  2548 => x"6000386c",
  2549 => x"00600000",
  2550 => x"0e006000",
  2551 => x"5d5c5b5e",
  2552 => x"4c711e0e",
  2553 => x"bfe6c6c3",
  2554 => x"eac6c34b",
  2555 => x"7478c048",
  2556 => x"c6e2c21e",
  2557 => x"c3e2fd1e",
  2558 => x"9786c887",
  2559 => x"0299496b",
  2560 => x"c087c8c1",
  2561 => x"eac6c31e",
  2562 => x"ad744dbf",
  2563 => x"c487c702",
  2564 => x"78c048a6",
  2565 => x"a6c487c5",
  2566 => x"c478c148",
  2567 => x"49751e66",
  2568 => x"c887feec",
  2569 => x"49e0c086",
  2570 => x"c487efee",
  2571 => x"496a4aa3",
  2572 => x"f087f1ef",
  2573 => x"c6c387c7",
  2574 => x"c148bfea",
  2575 => x"eec6c380",
  2576 => x"9783cc58",
  2577 => x"0599496b",
  2578 => x"c387f8fe",
  2579 => x"4dbfeac6",
  2580 => x"03adb7c8",
  2581 => x"1ec087d9",
  2582 => x"eac6c31e",
  2583 => x"c0ec49bf",
  2584 => x"ef86c887",
  2585 => x"85c187d7",
  2586 => x"04adb7c8",
  2587 => x"c387e7ff",
  2588 => x"1ebfeac6",
  2589 => x"1ed8e2c2",
  2590 => x"87c0e0fd",
  2591 => x"4d268ef4",
  2592 => x"4b264c26",
  2593 => x"69484f26",
  2594 => x"696c6867",
  2595 => x"20746867",
  2596 => x"20776f72",
  2597 => x"000a6425",
  2598 => x"756e654d",
  2599 => x"73616820",
  2600 => x"20642520",
  2601 => x"73776f72",
  2602 => x"6143000a",
  2603 => x"61626c6c",
  2604 => x"25206b63",
  2605 => x"45000a78",
  2606 => x"7265746e",
  2607 => x"74656420",
  2608 => x"65746365",
  2609 => x"64252064",
  2610 => x"63202d20",
  2611 => x"65727275",
  2612 => x"6f72746e",
  2613 => x"64252077",
  2614 => x"711e000a",
  2615 => x"eac6c34a",
  2616 => x"eec6c35a",
  2617 => x"f2fb49bf",
  2618 => x"eac6c387",
  2619 => x"89c149bf",
  2620 => x"59f2c6c3",
  2621 => x"87e3fb71",
  2622 => x"c11e4f26",
  2623 => x"f0e849c0",
  2624 => x"fff1c287",
  2625 => x"2678c048",
  2626 => x"5b5e0e4f",
  2627 => x"4bc00e5c",
  2628 => x"49dac14c",
  2629 => x"7087e5e4",
  2630 => x"87c30298",
  2631 => x"c14bc0c2",
  2632 => x"d7e449d9",
  2633 => x"02987087",
  2634 => x"c0c187c3",
  2635 => x"49d4c2b3",
  2636 => x"7087c9e4",
  2637 => x"87c20298",
  2638 => x"d1c2b3d0",
  2639 => x"87fce349",
  2640 => x"c3029870",
  2641 => x"b3e0c087",
  2642 => x"e349f5c3",
  2643 => x"987087ee",
  2644 => x"c887c202",
  2645 => x"49f2c34b",
  2646 => x"7087e1e3",
  2647 => x"87c20298",
  2648 => x"ebc3b3c4",
  2649 => x"87d4e349",
  2650 => x"c2029870",
  2651 => x"c3b3c287",
  2652 => x"c7e349f4",
  2653 => x"02987087",
  2654 => x"b3c187c2",
  2655 => x"e249d8c1",
  2656 => x"987087fa",
  2657 => x"c287c302",
  2658 => x"49d24cc0",
  2659 => x"7087ede2",
  2660 => x"87c30298",
  2661 => x"d4b4c0c1",
  2662 => x"87e0e249",
  2663 => x"c2029870",
  2664 => x"d1b4d087",
  2665 => x"87d4e249",
  2666 => x"c3029870",
  2667 => x"b4e0c087",
  2668 => x"c7e249dd",
  2669 => x"02987087",
  2670 => x"4cc887c2",
  2671 => x"fbe149db",
  2672 => x"02987087",
  2673 => x"b4c487c2",
  2674 => x"efe149dc",
  2675 => x"02987087",
  2676 => x"b4c287c2",
  2677 => x"e149e3c0",
  2678 => x"987087e2",
  2679 => x"c187c202",
  2680 => x"c01e73b4",
  2681 => x"87fce349",
  2682 => x"49c11e74",
  2683 => x"f887f5e3",
  2684 => x"87ccfa8e",
  2685 => x"5c5b5e0e",
  2686 => x"86f00e5d",
  2687 => x"c048a6c8",
  2688 => x"c080c478",
  2689 => x"c380f878",
  2690 => x"78bfe6c6",
  2691 => x"bff2c6c3",
  2692 => x"e049c74c",
  2693 => x"497087e6",
  2694 => x"d70299c2",
  2695 => x"fff1c287",
  2696 => x"bac14abf",
  2697 => x"5ac3f2c2",
  2698 => x"49a2c0c1",
  2699 => x"cc87c2e4",
  2700 => x"78c148a6",
  2701 => x"bffff1c2",
  2702 => x"fb87d905",
  2703 => x"fdc387cb",
  2704 => x"f7dfff49",
  2705 => x"49fac387",
  2706 => x"87f0dfff",
  2707 => x"bffff1c2",
  2708 => x"87e6c848",
  2709 => x"ff49f5c3",
  2710 => x"7087e1df",
  2711 => x"0299c249",
  2712 => x"c387ecc0",
  2713 => x"02bfeec6",
  2714 => x"c14887c9",
  2715 => x"f2c6c388",
  2716 => x"c387d758",
  2717 => x"49bfeac6",
  2718 => x"66c491cc",
  2719 => x"7ea1c881",
  2720 => x"c502bf6e",
  2721 => x"49ff4b87",
  2722 => x"a6cc0f73",
  2723 => x"c378c148",
  2724 => x"deff49f2",
  2725 => x"497087e6",
  2726 => x"c00299c2",
  2727 => x"a6cc87fb",
  2728 => x"eac6c348",
  2729 => x"66cc78bf",
  2730 => x"c389c149",
  2731 => x"7ebfeec6",
  2732 => x"06a9b76e",
  2733 => x"c14887c9",
  2734 => x"f2c6c380",
  2735 => x"cc87d558",
  2736 => x"91cc4966",
  2737 => x"c88166c4",
  2738 => x"bf6e7ea1",
  2739 => x"4b87c502",
  2740 => x"0f7349fe",
  2741 => x"c148a6cc",
  2742 => x"49fdc378",
  2743 => x"87dcddff",
  2744 => x"99c24970",
  2745 => x"87ecc002",
  2746 => x"bfeec6c3",
  2747 => x"c387c802",
  2748 => x"c048eec6",
  2749 => x"c387d878",
  2750 => x"49bfeac6",
  2751 => x"66c491cc",
  2752 => x"7ea1c881",
  2753 => x"c002bf6e",
  2754 => x"fd4b87c5",
  2755 => x"cc0f7349",
  2756 => x"78c148a6",
  2757 => x"ff49fac3",
  2758 => x"7087e1dc",
  2759 => x"0299c249",
  2760 => x"cc87ffc0",
  2761 => x"c6c348a6",
  2762 => x"cc78bfea",
  2763 => x"88c14866",
  2764 => x"c358a6c4",
  2765 => x"48bfeec6",
  2766 => x"03a8b76e",
  2767 => x"c387c8c0",
  2768 => x"6e48eec6",
  2769 => x"cc87d678",
  2770 => x"91cc4966",
  2771 => x"c88166c4",
  2772 => x"bf6e7ea1",
  2773 => x"87c5c002",
  2774 => x"7349fc4b",
  2775 => x"48a6cc0f",
  2776 => x"c6c378c1",
  2777 => x"c04bbfee",
  2778 => x"c006abb7",
  2779 => x"8bc187c9",
  2780 => x"01abb7c0",
  2781 => x"c187f7ff",
  2782 => x"daff49da",
  2783 => x"497087fe",
  2784 => x"739bc24b",
  2785 => x"f1c2029b",
  2786 => x"e6c6c387",
  2787 => x"c6c34dbf",
  2788 => x"731ebfee",
  2789 => x"f7e2c21e",
  2790 => x"dfd3fd1e",
  2791 => x"c386cc87",
  2792 => x"4bbfeec6",
  2793 => x"06abb7c0",
  2794 => x"cc87cbc0",
  2795 => x"c08bc185",
  2796 => x"ff01abb7",
  2797 => x"6d9787f5",
  2798 => x"028ac14a",
  2799 => x"8a87f5c0",
  2800 => x"87d5c002",
  2801 => x"cbc1028a",
  2802 => x"c1058a87",
  2803 => x"a5c887ec",
  2804 => x"f4496a4a",
  2805 => x"e1c187c4",
  2806 => x"4ba5c887",
  2807 => x"e2c21e6b",
  2808 => x"d2fd1eea",
  2809 => x"86c887d6",
  2810 => x"c6c34b6b",
  2811 => x"7349bfee",
  2812 => x"87c6c10f",
  2813 => x"c149a5c8",
  2814 => x"70306948",
  2815 => x"e2c6c349",
  2816 => x"b87148bf",
  2817 => x"58e6c6c3",
  2818 => x"c148a6cc",
  2819 => x"c180fc78",
  2820 => x"87e6c078",
  2821 => x"cb49a5c8",
  2822 => x"976e7ea5",
  2823 => x"a2c14abf",
  2824 => x"4969974b",
  2825 => x"c004abb7",
  2826 => x"4bc087c2",
  2827 => x"7b970b6e",
  2828 => x"48a6cc0b",
  2829 => x"80fc78c1",
  2830 => x"9c7478c1",
  2831 => x"87e9c002",
  2832 => x"e4c0026c",
  2833 => x"ff496c87",
  2834 => x"7087f1d7",
  2835 => x"0299c149",
  2836 => x"c487cbc0",
  2837 => x"c6c34ba4",
  2838 => x"6b49bfee",
  2839 => x"84c80f4b",
  2840 => x"87c5c002",
  2841 => x"dcff056c",
  2842 => x"0266cc87",
  2843 => x"c387c8c0",
  2844 => x"49bfeec6",
  2845 => x"c887e4ed",
  2846 => x"8ef04866",
  2847 => x"0087ffef",
  2848 => x"b1000000",
  2849 => x"b100001f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
