library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0c1c387",
    12 => x"86c0d04e",
    13 => x"49c0c1c3",
    14 => x"48ccecc2",
    15 => x"0389d089",
    16 => x"404040c0",
    17 => x"d087f640",
    18 => x"50c00581",
    19 => x"f90589c1",
    20 => x"ccecc287",
    21 => x"c8ecc24d",
    22 => x"02ad744c",
    23 => x"0f2487c4",
    24 => x"f3c187f7",
    25 => x"ecc287d5",
    26 => x"ecc24dcc",
    27 => x"ad744ccc",
    28 => x"c487c602",
    29 => x"f50f6c8c",
    30 => x"87fd0087",
    31 => x"5c5b5e0e",
    32 => x"86f00e5d",
    33 => x"a6c44cc0",
    34 => x"c078c048",
    35 => x"c04ba6e4",
    36 => x"484966e0",
    37 => x"e4c080c1",
    38 => x"481158a6",
    39 => x"7058a6c4",
    40 => x"f6c30298",
    41 => x"0266c487",
    42 => x"c487c6c3",
    43 => x"78c048a6",
    44 => x"f0c04a6e",
    45 => x"dac2028a",
    46 => x"8af3c087",
    47 => x"87dbc202",
    48 => x"dc028ac1",
    49 => x"028ac887",
    50 => x"c487c8c2",
    51 => x"87d1028a",
    52 => x"c1028ac3",
    53 => x"8ac287eb",
    54 => x"c387c602",
    55 => x"c9c2058a",
    56 => x"7383c487",
    57 => x"6989c449",
    58 => x"c1026e7e",
    59 => x"a6c887c8",
    60 => x"c478c048",
    61 => x"cc78c080",
    62 => x"4a6e4d66",
    63 => x"cf2ab7dc",
    64 => x"c4486e9a",
    65 => x"7258a630",
    66 => x"87c5029a",
    67 => x"c148a6c8",
    68 => x"06aac978",
    69 => x"f7c087c5",
    70 => x"c087c382",
    71 => x"66c882f0",
    72 => x"7287c702",
    73 => x"87f3c249",
    74 => x"85c184c1",
    75 => x"04adb7c8",
    76 => x"c187c7ff",
    77 => x"f0c087cf",
    78 => x"87dfc249",
    79 => x"c4c184c1",
    80 => x"7383c487",
    81 => x"6a8ac44a",
    82 => x"87dbc149",
    83 => x"4ca44970",
    84 => x"c487f2c0",
    85 => x"78c148a6",
    86 => x"c487eac0",
    87 => x"c44a7383",
    88 => x"c1496a8a",
    89 => x"84c187f5",
    90 => x"496e87db",
    91 => x"d487ecc1",
    92 => x"c0486e87",
    93 => x"c705a8e5",
    94 => x"48a6c487",
    95 => x"87c578c1",
    96 => x"d6c1496e",
    97 => x"66e0c087",
    98 => x"80c14849",
    99 => x"58a6e4c0",
   100 => x"a6c44811",
   101 => x"05987058",
   102 => x"7487cafc",
   103 => x"268ef048",
   104 => x"264c264d",
   105 => x"0e4f264b",
   106 => x"0e5c5b5e",
   107 => x"4cc04b71",
   108 => x"029a4a13",
   109 => x"497287cd",
   110 => x"c187e0c0",
   111 => x"9a4a1384",
   112 => x"7487f305",
   113 => x"264c2648",
   114 => x"1e4f264b",
   115 => x"73814873",
   116 => x"87c502a9",
   117 => x"f6055312",
   118 => x"1e4f2687",
   119 => x"4ac0ff1e",
   120 => x"c0c4486a",
   121 => x"58a6c498",
   122 => x"f3029870",
   123 => x"487a7187",
   124 => x"1e4f2626",
   125 => x"d4ff1e73",
   126 => x"7bffc34b",
   127 => x"ffc34a6b",
   128 => x"c8496b7b",
   129 => x"c3b17232",
   130 => x"4a6b7bff",
   131 => x"b27131c8",
   132 => x"6b7bffc3",
   133 => x"7232c849",
   134 => x"c44871b1",
   135 => x"264d2687",
   136 => x"264b264c",
   137 => x"5b5e0e4f",
   138 => x"710e5d5c",
   139 => x"4cd4ff4a",
   140 => x"ffc34872",
   141 => x"c27c7098",
   142 => x"05bfccec",
   143 => x"66d087c8",
   144 => x"d430c948",
   145 => x"66d058a6",
   146 => x"7129d849",
   147 => x"98ffc348",
   148 => x"66d07c70",
   149 => x"7129d049",
   150 => x"98ffc348",
   151 => x"66d07c70",
   152 => x"7129c849",
   153 => x"98ffc348",
   154 => x"66d07c70",
   155 => x"98ffc348",
   156 => x"49727c70",
   157 => x"487129d0",
   158 => x"7098ffc3",
   159 => x"c94b6c7c",
   160 => x"c34dfff0",
   161 => x"d005abff",
   162 => x"7cffc387",
   163 => x"8dc14b6c",
   164 => x"c387c602",
   165 => x"f002abff",
   166 => x"fd487387",
   167 => x"c01e87ff",
   168 => x"48d4ff49",
   169 => x"c178ffc3",
   170 => x"b7c8c381",
   171 => x"87f104a9",
   172 => x"731e4f26",
   173 => x"c487e71e",
   174 => x"c04bdff8",
   175 => x"f0ffc01e",
   176 => x"fd49f7c1",
   177 => x"86c487df",
   178 => x"c005a8c1",
   179 => x"d4ff87ea",
   180 => x"78ffc348",
   181 => x"c0c0c0c1",
   182 => x"c01ec0c0",
   183 => x"e9c1f0e1",
   184 => x"87c1fd49",
   185 => x"987086c4",
   186 => x"ff87ca05",
   187 => x"ffc348d4",
   188 => x"cb48c178",
   189 => x"87e6fe87",
   190 => x"fe058bc1",
   191 => x"48c087fd",
   192 => x"1e87defc",
   193 => x"d4ff1e73",
   194 => x"78ffc348",
   195 => x"fa49fecc",
   196 => x"4bd387d5",
   197 => x"ffc01ec0",
   198 => x"49c1c1f0",
   199 => x"c487c6fc",
   200 => x"05987086",
   201 => x"d4ff87ca",
   202 => x"78ffc348",
   203 => x"87cb48c1",
   204 => x"c187ebfd",
   205 => x"dbff058b",
   206 => x"fb48c087",
   207 => x"4d4387e3",
   208 => x"4d430044",
   209 => x"20383544",
   210 => x"200a6425",
   211 => x"4d430020",
   212 => x"5f383544",
   213 => x"64252032",
   214 => x"0020200a",
   215 => x"35444d43",
   216 => x"64252038",
   217 => x"0020200a",
   218 => x"43484453",
   219 => x"696e4920",
   220 => x"6c616974",
   221 => x"74617a69",
   222 => x"206e6f69",
   223 => x"6f727265",
   224 => x"000a2172",
   225 => x"5f646d63",
   226 => x"38444d43",
   227 => x"73657220",
   228 => x"736e6f70",
   229 => x"25203a65",
   230 => x"49000a64",
   231 => x"00525245",
   232 => x"00495053",
   233 => x"63204453",
   234 => x"20647261",
   235 => x"657a6973",
   236 => x"20736920",
   237 => x"000a6425",
   238 => x"74697257",
   239 => x"61662065",
   240 => x"64656c69",
   241 => x"5f63000a",
   242 => x"657a6973",
   243 => x"6c756d5f",
   244 => x"25203a74",
   245 => x"72202c64",
   246 => x"5f646165",
   247 => x"6c5f6c62",
   248 => x"203a6e65",
   249 => x"202c6425",
   250 => x"7a697363",
   251 => x"25203a65",
   252 => x"4d000a64",
   253 => x"20746c75",
   254 => x"000a6425",
   255 => x"62206425",
   256 => x"6b636f6c",
   257 => x"666f2073",
   258 => x"7a697320",
   259 => x"64252065",
   260 => x"6425000a",
   261 => x"6f6c6220",
   262 => x"20736b63",
   263 => x"3520666f",
   264 => x"62203231",
   265 => x"73657479",
   266 => x"5e0e000a",
   267 => x"0e5d5c5b",
   268 => x"f94dd4ff",
   269 => x"eac687e8",
   270 => x"f0e1c01e",
   271 => x"f749c8c1",
   272 => x"4b7087e3",
   273 => x"1ec4ce1e",
   274 => x"cc87f1f0",
   275 => x"02abc186",
   276 => x"eefa87c8",
   277 => x"c248c087",
   278 => x"d6f687ca",
   279 => x"cf497087",
   280 => x"c699ffff",
   281 => x"c802a9ea",
   282 => x"87d7fa87",
   283 => x"f3c148c0",
   284 => x"7dffc387",
   285 => x"f84cf1c0",
   286 => x"987087f8",
   287 => x"87cbc102",
   288 => x"ffc01ec0",
   289 => x"49fac1f0",
   290 => x"c487daf6",
   291 => x"9b4b7086",
   292 => x"87edc005",
   293 => x"1ec2cd1e",
   294 => x"c387e1ef",
   295 => x"4b6d7dff",
   296 => x"1ececd1e",
   297 => x"d087d5ef",
   298 => x"7dffc386",
   299 => x"737d7d7d",
   300 => x"99c0c149",
   301 => x"c187c502",
   302 => x"87e8c048",
   303 => x"e3c048c0",
   304 => x"cd1e7387",
   305 => x"f3ee1edc",
   306 => x"c286c887",
   307 => x"87cc05ac",
   308 => x"ee1ee8cd",
   309 => x"86c487e6",
   310 => x"87c848c0",
   311 => x"fe058cc1",
   312 => x"48c087d5",
   313 => x"0e87f6f4",
   314 => x"5d5c5b5e",
   315 => x"d0ff1e0e",
   316 => x"c0c0c84d",
   317 => x"ccecc24b",
   318 => x"ce78c148",
   319 => x"e6f249e0",
   320 => x"6d4cc787",
   321 => x"c4987348",
   322 => x"987058a6",
   323 => x"6d87cc02",
   324 => x"c4987348",
   325 => x"987058a6",
   326 => x"c287f405",
   327 => x"87fef57d",
   328 => x"9873486d",
   329 => x"7058a6c4",
   330 => x"87cc0298",
   331 => x"9873486d",
   332 => x"7058a6c4",
   333 => x"87f40598",
   334 => x"1ec07dc3",
   335 => x"c1d0e5c0",
   336 => x"e0f349c0",
   337 => x"c186c487",
   338 => x"87c105a8",
   339 => x"05acc24c",
   340 => x"dbce87cb",
   341 => x"87cff149",
   342 => x"d8c148c0",
   343 => x"058cc187",
   344 => x"fb87e0fe",
   345 => x"ecc287c4",
   346 => x"987058d0",
   347 => x"c187cd05",
   348 => x"f0ffc01e",
   349 => x"f249d0c1",
   350 => x"86c487eb",
   351 => x"c348d4ff",
   352 => x"e7c578ff",
   353 => x"d4ecc287",
   354 => x"ce1e7058",
   355 => x"ebeb1ee4",
   356 => x"6d86c887",
   357 => x"c4987348",
   358 => x"987058a6",
   359 => x"6d87cc02",
   360 => x"c4987348",
   361 => x"987058a6",
   362 => x"c287f405",
   363 => x"48d4ff7d",
   364 => x"c178ffc3",
   365 => x"e4f12648",
   366 => x"5b5e0e87",
   367 => x"1e0e5d5c",
   368 => x"4bc0c0c8",
   369 => x"eec54cc0",
   370 => x"c44adfcd",
   371 => x"d4ff5ca6",
   372 => x"7cffc34c",
   373 => x"fec3486c",
   374 => x"c0c205a8",
   375 => x"05997187",
   376 => x"ff87e2c0",
   377 => x"7348bfd0",
   378 => x"58a6c498",
   379 => x"ce029870",
   380 => x"bfd0ff87",
   381 => x"c4987348",
   382 => x"987058a6",
   383 => x"ff87f205",
   384 => x"d1c448d0",
   385 => x"4866d478",
   386 => x"06a8b7c0",
   387 => x"c387e0c0",
   388 => x"4a6c7cff",
   389 => x"c7029971",
   390 => x"970a7187",
   391 => x"81c10a7a",
   392 => x"c14866d4",
   393 => x"58a6d888",
   394 => x"01a8b7c0",
   395 => x"c387e0ff",
   396 => x"717c7cff",
   397 => x"e1c00599",
   398 => x"bfd0ff87",
   399 => x"c4987348",
   400 => x"987058a6",
   401 => x"ff87ce02",
   402 => x"7348bfd0",
   403 => x"58a6c498",
   404 => x"f2059870",
   405 => x"48d0ff87",
   406 => x"4ac178d0",
   407 => x"058ac17e",
   408 => x"6e87eefd",
   409 => x"f4ee2648",
   410 => x"5b5e0e87",
   411 => x"711e0e5c",
   412 => x"c0c0c84a",
   413 => x"ff4cc04b",
   414 => x"ffc348d4",
   415 => x"bfd0ff78",
   416 => x"c4987348",
   417 => x"987058a6",
   418 => x"ff87ce02",
   419 => x"7348bfd0",
   420 => x"58a6c498",
   421 => x"f2059870",
   422 => x"48d0ff87",
   423 => x"ff78c3c4",
   424 => x"ffc348d4",
   425 => x"c01e7278",
   426 => x"d1c1f0ff",
   427 => x"87f5ed49",
   428 => x"987086c4",
   429 => x"87eec005",
   430 => x"d41ec0c8",
   431 => x"f8fb4966",
   432 => x"7086c487",
   433 => x"bfd0ff4c",
   434 => x"c4987348",
   435 => x"987058a6",
   436 => x"ff87ce02",
   437 => x"7348bfd0",
   438 => x"58a6c498",
   439 => x"f2059870",
   440 => x"48d0ff87",
   441 => x"487478c2",
   442 => x"87f3ec26",
   443 => x"5c5b5e0e",
   444 => x"c01e0e5d",
   445 => x"f0ffc01e",
   446 => x"ec49c9c1",
   447 => x"1ed287e7",
   448 => x"49daecc2",
   449 => x"c887f2fa",
   450 => x"c14dc086",
   451 => x"adb7d285",
   452 => x"c287f804",
   453 => x"bf97daec",
   454 => x"99c0c349",
   455 => x"05a9c0c1",
   456 => x"c287e7c0",
   457 => x"bf97e1ec",
   458 => x"c231d049",
   459 => x"bf97e2ec",
   460 => x"7232c84a",
   461 => x"e3ecc2b1",
   462 => x"b14abf97",
   463 => x"ffcf4d71",
   464 => x"c19dffff",
   465 => x"c235ca85",
   466 => x"ecc287de",
   467 => x"4bbf97e3",
   468 => x"9bc633c1",
   469 => x"97e4ecc2",
   470 => x"b7c749bf",
   471 => x"c2b37129",
   472 => x"bf97dfec",
   473 => x"98cf4849",
   474 => x"c258a6c4",
   475 => x"bf97e0ec",
   476 => x"ca9cc34c",
   477 => x"e1ecc234",
   478 => x"c249bf97",
   479 => x"c2b47131",
   480 => x"bf97e2ec",
   481 => x"99c0c349",
   482 => x"7129b7c6",
   483 => x"701e74b4",
   484 => x"cf1e731e",
   485 => x"e3e31ec6",
   486 => x"c183c287",
   487 => x"70307348",
   488 => x"f3cf1e4b",
   489 => x"87d4e31e",
   490 => x"66d848c1",
   491 => x"58a6dc30",
   492 => x"4d49a4c1",
   493 => x"1e709573",
   494 => x"fccf1e75",
   495 => x"87fce21e",
   496 => x"6e86e4c0",
   497 => x"b7c0c848",
   498 => x"87d206a8",
   499 => x"486e35c1",
   500 => x"c428b7c1",
   501 => x"c0c858a6",
   502 => x"ff01a8b7",
   503 => x"1e7587ee",
   504 => x"e21ed2d0",
   505 => x"86c887d6",
   506 => x"e8264875",
   507 => x"5e0e87ef",
   508 => x"710e5c5b",
   509 => x"d04cc04b",
   510 => x"b7c04866",
   511 => x"e3c006a8",
   512 => x"cc4a1387",
   513 => x"49bf9766",
   514 => x"c14866cc",
   515 => x"58a6d080",
   516 => x"02aab771",
   517 => x"48c187c4",
   518 => x"84c187cc",
   519 => x"acb766d0",
   520 => x"87ddff04",
   521 => x"87c248c0",
   522 => x"4c264d26",
   523 => x"4f264b26",
   524 => x"5c5b5e0e",
   525 => x"f5c20e5d",
   526 => x"78c048c0",
   527 => x"49ddefc0",
   528 => x"c287e4e5",
   529 => x"c01ef8ec",
   530 => x"87ddf849",
   531 => x"987086c4",
   532 => x"c087cc05",
   533 => x"e549c9ec",
   534 => x"48c087cd",
   535 => x"c087e7ca",
   536 => x"e549eaef",
   537 => x"4bc087c1",
   538 => x"48f8f9c2",
   539 => x"1ec878c1",
   540 => x"1ec1f0c0",
   541 => x"49eeedc2",
   542 => x"c887f3fd",
   543 => x"05987086",
   544 => x"f9c287c6",
   545 => x"78c048f8",
   546 => x"f0c01ec8",
   547 => x"eec21eca",
   548 => x"d9fd49ca",
   549 => x"7086c887",
   550 => x"87c60598",
   551 => x"48f8f9c2",
   552 => x"f9c278c0",
   553 => x"c01ebff8",
   554 => x"ff1ed3f0",
   555 => x"c887cddf",
   556 => x"f8f9c286",
   557 => x"f7c102bf",
   558 => x"f6f4c287",
   559 => x"1e49bf9f",
   560 => x"49f6f4c2",
   561 => x"a0c2f848",
   562 => x"d01e7189",
   563 => x"1ec0c81e",
   564 => x"1efbecc0",
   565 => x"87e4deff",
   566 => x"f3c286d4",
   567 => x"c24bbffe",
   568 => x"bf9ff6f4",
   569 => x"ead6c54a",
   570 => x"c8c005aa",
   571 => x"fef3c287",
   572 => x"d4c04bbf",
   573 => x"d5e9ca87",
   574 => x"ccc002aa",
   575 => x"ddecc087",
   576 => x"87e3e249",
   577 => x"fdc748c0",
   578 => x"c01e7387",
   579 => x"ff1ef8ed",
   580 => x"c287e9dd",
   581 => x"731ef8ec",
   582 => x"87cdf549",
   583 => x"987086cc",
   584 => x"87c5c005",
   585 => x"ddc748c0",
   586 => x"d0eec087",
   587 => x"87f7e149",
   588 => x"1ee6f0c0",
   589 => x"87c4ddff",
   590 => x"f0c01ec8",
   591 => x"eec21efe",
   592 => x"e9fa49ca",
   593 => x"7086cc87",
   594 => x"c9c00598",
   595 => x"c0f5c287",
   596 => x"c078c148",
   597 => x"1ec887e4",
   598 => x"1ec7f1c0",
   599 => x"49eeedc2",
   600 => x"c887cbfa",
   601 => x"02987086",
   602 => x"c087cfc0",
   603 => x"ff1ef7ee",
   604 => x"c487c9dc",
   605 => x"c648c086",
   606 => x"f4c287cc",
   607 => x"49bf97f6",
   608 => x"05a9d5c1",
   609 => x"c287cdc0",
   610 => x"bf97f7f4",
   611 => x"a9eac249",
   612 => x"87c5c002",
   613 => x"edc548c0",
   614 => x"f8ecc287",
   615 => x"c34cbf97",
   616 => x"c002ace9",
   617 => x"ebc387cc",
   618 => x"c5c002ac",
   619 => x"c548c087",
   620 => x"edc287d4",
   621 => x"49bf97c3",
   622 => x"ccc00599",
   623 => x"c4edc287",
   624 => x"c249bf97",
   625 => x"c5c002a9",
   626 => x"c448c087",
   627 => x"edc287f8",
   628 => x"48bf97c5",
   629 => x"58fcf4c2",
   630 => x"c14a4970",
   631 => x"c0f5c28a",
   632 => x"711e725a",
   633 => x"d0f1c01e",
   634 => x"cfdaff1e",
   635 => x"c286cc87",
   636 => x"bf97c6ed",
   637 => x"c2817349",
   638 => x"bf97c7ed",
   639 => x"35c84d4a",
   640 => x"f9c28571",
   641 => x"edc25dd8",
   642 => x"48bf97c8",
   643 => x"58ecf9c2",
   644 => x"bfc0f5c2",
   645 => x"87dcc202",
   646 => x"efc01ec8",
   647 => x"eec21ed4",
   648 => x"c9f749ca",
   649 => x"7086c887",
   650 => x"c5c00298",
   651 => x"c348c087",
   652 => x"f4c287d4",
   653 => x"484abff8",
   654 => x"f5c230c4",
   655 => x"f9c258c8",
   656 => x"edc25ae8",
   657 => x"49bf97dd",
   658 => x"edc231c8",
   659 => x"4bbf97dc",
   660 => x"edc249a1",
   661 => x"4bbf97de",
   662 => x"a17333d0",
   663 => x"dfedc249",
   664 => x"d84bbf97",
   665 => x"49a17333",
   666 => x"59f0f9c2",
   667 => x"bfe8f9c2",
   668 => x"d4f9c291",
   669 => x"f9c281bf",
   670 => x"edc259dc",
   671 => x"4bbf97e5",
   672 => x"edc233c8",
   673 => x"4cbf97e4",
   674 => x"edc24ba3",
   675 => x"4cbf97e6",
   676 => x"a37434d0",
   677 => x"e7edc24b",
   678 => x"cf4cbf97",
   679 => x"7434d89c",
   680 => x"f9c24ba3",
   681 => x"8bc25be0",
   682 => x"f9c29273",
   683 => x"a17248e0",
   684 => x"87cbc178",
   685 => x"97caedc2",
   686 => x"31c849bf",
   687 => x"97c9edc2",
   688 => x"49a14abf",
   689 => x"59c8f5c2",
   690 => x"ffc731c5",
   691 => x"c229c981",
   692 => x"c259e8f9",
   693 => x"bf97cfed",
   694 => x"c232c84a",
   695 => x"bf97ceed",
   696 => x"c24aa24b",
   697 => x"c25af0f9",
   698 => x"92bfe8f9",
   699 => x"f9c28275",
   700 => x"f9c25ae4",
   701 => x"78c048dc",
   702 => x"48d8f9c2",
   703 => x"c078a172",
   704 => x"87e3cd49",
   705 => x"dff448c1",
   706 => x"61655287",
   707 => x"666f2064",
   708 => x"52424d20",
   709 => x"69616620",
   710 => x"0a64656c",
   711 => x"206f4e00",
   712 => x"74726170",
   713 => x"6f697469",
   714 => x"6973206e",
   715 => x"74616e67",
   716 => x"20657275",
   717 => x"6e756f66",
   718 => x"4d000a64",
   719 => x"69735242",
   720 => x"203a657a",
   721 => x"202c6425",
   722 => x"74726170",
   723 => x"6f697469",
   724 => x"7a69736e",
   725 => x"25203a65",
   726 => x"6f202c64",
   727 => x"65736666",
   728 => x"666f2074",
   729 => x"67697320",
   730 => x"6425203a",
   731 => x"6973202c",
   732 => x"78302067",
   733 => x"000a7825",
   734 => x"64616552",
   735 => x"20676e69",
   736 => x"746f6f62",
   737 => x"63657320",
   738 => x"20726f74",
   739 => x"000a6425",
   740 => x"64616552",
   741 => x"6f6f6220",
   742 => x"65732074",
   743 => x"726f7463",
   744 => x"6f726620",
   745 => x"6966206d",
   746 => x"20747372",
   747 => x"74726170",
   748 => x"6f697469",
   749 => x"55000a6e",
   750 => x"7075736e",
   751 => x"74726f70",
   752 => x"70206465",
   753 => x"69747261",
   754 => x"6e6f6974",
   755 => x"70797420",
   756 => x"000d2165",
   757 => x"33544146",
   758 => x"20202032",
   759 => x"61655200",
   760 => x"676e6964",
   761 => x"52424d20",
   762 => x"424d000a",
   763 => x"75732052",
   764 => x"73656363",
   765 => x"6c756673",
   766 => x"7220796c",
   767 => x"0a646165",
   768 => x"54414600",
   769 => x"20203631",
   770 => x"41460020",
   771 => x"20323354",
   772 => x"50002020",
   773 => x"69747261",
   774 => x"6e6f6974",
   775 => x"6e756f63",
   776 => x"64252074",
   777 => x"7548000a",
   778 => x"6e69746e",
   779 => x"6f662067",
   780 => x"69662072",
   781 => x"7973656c",
   782 => x"6d657473",
   783 => x"4146000a",
   784 => x"20323354",
   785 => x"46002020",
   786 => x"36315441",
   787 => x"00202020",
   788 => x"73756c43",
   789 => x"20726574",
   790 => x"657a6973",
   791 => x"6425203a",
   792 => x"6c43202c",
   793 => x"65747375",
   794 => x"616d2072",
   795 => x"202c6b73",
   796 => x"000a6425",
   797 => x"6e65704f",
   798 => x"66206465",
   799 => x"2c656c69",
   800 => x"616f6c20",
   801 => x"676e6964",
   802 => x"0a2e2e2e",
   803 => x"6e614300",
   804 => x"6f207427",
   805 => x"206e6570",
   806 => x"000a7325",
   807 => x"5c5b5e0e",
   808 => x"4a710e5d",
   809 => x"bfc0f5c2",
   810 => x"7287cc02",
   811 => x"2bb7c74b",
   812 => x"ffc14d72",
   813 => x"7287ca9d",
   814 => x"2bb7c84b",
   815 => x"ffc34d72",
   816 => x"f8ecc29d",
   817 => x"d4f9c21e",
   818 => x"817349bf",
   819 => x"87d9e671",
   820 => x"987086c4",
   821 => x"c087c505",
   822 => x"87e6c048",
   823 => x"bfc0f5c2",
   824 => x"7587d202",
   825 => x"c291c449",
   826 => x"6981f8ec",
   827 => x"ffffcf4c",
   828 => x"cb9cffff",
   829 => x"c2497587",
   830 => x"f8ecc291",
   831 => x"4c699f81",
   832 => x"e3ec4874",
   833 => x"5b5e0e87",
   834 => x"f40e5d5c",
   835 => x"c04c7186",
   836 => x"f0f9c24b",
   837 => x"a6c47ebf",
   838 => x"f4f9c248",
   839 => x"a6c878bf",
   840 => x"c278c048",
   841 => x"48bfc4f5",
   842 => x"c206a8c0",
   843 => x"66c887e3",
   844 => x"0599cf49",
   845 => x"ecc287d8",
   846 => x"66c81ef8",
   847 => x"80c14849",
   848 => x"e458a6cc",
   849 => x"86c487e3",
   850 => x"4bf8ecc2",
   851 => x"e0c087c3",
   852 => x"4a6b9783",
   853 => x"e7c1029a",
   854 => x"aae5c387",
   855 => x"87e0c102",
   856 => x"9749a3cb",
   857 => x"99d84969",
   858 => x"87d4c105",
   859 => x"d0ff4973",
   860 => x"1ecb87f5",
   861 => x"1e66e0c0",
   862 => x"f1e94973",
   863 => x"7086c887",
   864 => x"fbc00598",
   865 => x"4aa3dc87",
   866 => x"6a49a4c4",
   867 => x"49a3da79",
   868 => x"9f4da4c8",
   869 => x"c27d4869",
   870 => x"02bfc0f5",
   871 => x"a3d487d3",
   872 => x"49699f49",
   873 => x"99ffffc0",
   874 => x"30d04871",
   875 => x"c258a6c4",
   876 => x"6e7ec087",
   877 => x"70806d48",
   878 => x"c17cc07d",
   879 => x"87c5c148",
   880 => x"c14866c8",
   881 => x"58a6cc80",
   882 => x"bfc4f5c2",
   883 => x"ddfd04a8",
   884 => x"c0f5c287",
   885 => x"eac002bf",
   886 => x"fa496e87",
   887 => x"a6c487fe",
   888 => x"cf497058",
   889 => x"f8ffffff",
   890 => x"d602a999",
   891 => x"c2497087",
   892 => x"f8f4c289",
   893 => x"f9c291bf",
   894 => x"7148bfd8",
   895 => x"58a6c880",
   896 => x"c087dbfc",
   897 => x"e88ef448",
   898 => x"731e87de",
   899 => x"6a4a711e",
   900 => x"7181c149",
   901 => x"fcf4c27a",
   902 => x"cb0599bf",
   903 => x"4ba2c887",
   904 => x"f7f9496b",
   905 => x"7b497087",
   906 => x"ffe748c1",
   907 => x"1e731e87",
   908 => x"f9c24b71",
   909 => x"c849bfd8",
   910 => x"4a6a4aa3",
   911 => x"f4c28ac2",
   912 => x"7292bff8",
   913 => x"f4c249a1",
   914 => x"6b4abffc",
   915 => x"49a1729a",
   916 => x"711e66c8",
   917 => x"c487d2e0",
   918 => x"05987086",
   919 => x"48c087c4",
   920 => x"48c187c2",
   921 => x"0e87c5e7",
   922 => x"0e5c5b5e",
   923 => x"4bc04a71",
   924 => x"c0029a72",
   925 => x"a2da87e0",
   926 => x"4b699f49",
   927 => x"bfc0f5c2",
   928 => x"d487cf02",
   929 => x"699f49a2",
   930 => x"ffc04c49",
   931 => x"34d09cff",
   932 => x"4cc087c2",
   933 => x"9b73b374",
   934 => x"4a87df02",
   935 => x"f4c28ac2",
   936 => x"9249bff8",
   937 => x"bfd8f9c2",
   938 => x"c2807248",
   939 => x"7158f8f9",
   940 => x"c230c448",
   941 => x"c058c8f5",
   942 => x"f9c287e9",
   943 => x"c24bbfdc",
   944 => x"c248f4f9",
   945 => x"78bfe0f9",
   946 => x"bfc0f5c2",
   947 => x"c287c902",
   948 => x"49bff8f4",
   949 => x"87c731c4",
   950 => x"bfe4f9c2",
   951 => x"c231c449",
   952 => x"c259c8f5",
   953 => x"e55bf4f9",
   954 => x"5e0e87c0",
   955 => x"0e5d5c5b",
   956 => x"9a4a711e",
   957 => x"c287de02",
   958 => x"c048f4ec",
   959 => x"ececc278",
   960 => x"f4f9c248",
   961 => x"ecc278bf",
   962 => x"f9c248f0",
   963 => x"c178bff0",
   964 => x"c048e2c2",
   965 => x"c4f5c278",
   966 => x"ecc249bf",
   967 => x"714abff4",
   968 => x"fec303aa",
   969 => x"cf497287",
   970 => x"e1c00599",
   971 => x"f8ecc287",
   972 => x"ececc21e",
   973 => x"ecc249bf",
   974 => x"a1c148ec",
   975 => x"dcff7178",
   976 => x"86c487e7",
   977 => x"48dec2c1",
   978 => x"78f8ecc2",
   979 => x"c2c187cc",
   980 => x"c048bfde",
   981 => x"c2c180e0",
   982 => x"ecc258e2",
   983 => x"c148bff4",
   984 => x"f8ecc280",
   985 => x"dec2c158",
   986 => x"a3cb4bbf",
   987 => x"cf4c1149",
   988 => x"ddc105ac",
   989 => x"109e2787",
   990 => x"97bf0000",
   991 => x"99df49bf",
   992 => x"91cd89c1",
   993 => x"81c8f5c2",
   994 => x"124aa3c1",
   995 => x"4aa3c351",
   996 => x"a3c55112",
   997 => x"c751124a",
   998 => x"51124aa3",
   999 => x"124aa3c9",
  1000 => x"4aa3ce51",
  1001 => x"a3d05112",
  1002 => x"d251124a",
  1003 => x"51124aa3",
  1004 => x"124aa3d4",
  1005 => x"4aa3d651",
  1006 => x"a3d85112",
  1007 => x"dc51124a",
  1008 => x"51124aa3",
  1009 => x"124aa3de",
  1010 => x"e2c2c151",
  1011 => x"c178c148",
  1012 => x"497487c1",
  1013 => x"c00599c8",
  1014 => x"497487f3",
  1015 => x"d00599d0",
  1016 => x"0266d487",
  1017 => x"7387cac0",
  1018 => x"0f66d449",
  1019 => x"dc029870",
  1020 => x"e2c2c187",
  1021 => x"c6c005bf",
  1022 => x"c8f5c287",
  1023 => x"c150c048",
  1024 => x"c048e2c2",
  1025 => x"dec2c178",
  1026 => x"ccc248bf",
  1027 => x"e2c2c187",
  1028 => x"c278c048",
  1029 => x"49bfc4f5",
  1030 => x"bff4ecc2",
  1031 => x"04aa714a",
  1032 => x"c287c2fc",
  1033 => x"05bff4f9",
  1034 => x"c287c8c0",
  1035 => x"02bfc0f5",
  1036 => x"c287e4c1",
  1037 => x"49bff0ec",
  1038 => x"c287e1f1",
  1039 => x"7058f4ec",
  1040 => x"c0f5c24d",
  1041 => x"d7c002bf",
  1042 => x"cf497587",
  1043 => x"f8ffffff",
  1044 => x"c002a999",
  1045 => x"4cc087c5",
  1046 => x"c187d9c0",
  1047 => x"87d4c04c",
  1048 => x"ffcf4975",
  1049 => x"02a999f8",
  1050 => x"c087c5c0",
  1051 => x"87c2c07e",
  1052 => x"4c6e7ec1",
  1053 => x"c0059c74",
  1054 => x"497587dd",
  1055 => x"f4c289c2",
  1056 => x"c291bff8",
  1057 => x"48bfd8f9",
  1058 => x"ecc28071",
  1059 => x"ecc258f0",
  1060 => x"78c048f4",
  1061 => x"c087fef9",
  1062 => x"deff2648",
  1063 => x"000087ca",
  1064 => x"00000000",
  1065 => x"ff1e0000",
  1066 => x"ffc348d4",
  1067 => x"99496878",
  1068 => x"c087c602",
  1069 => x"ee05a9fb",
  1070 => x"26487187",
  1071 => x"5b5e0e4f",
  1072 => x"4a710e5c",
  1073 => x"d4ff4bc0",
  1074 => x"78ffc348",
  1075 => x"02994968",
  1076 => x"c087c1c1",
  1077 => x"c002a9ec",
  1078 => x"fbc087fa",
  1079 => x"f3c002a9",
  1080 => x"b766cc87",
  1081 => x"87cc03ab",
  1082 => x"c70266d0",
  1083 => x"97097287",
  1084 => x"82c10979",
  1085 => x"c2029971",
  1086 => x"ff83c187",
  1087 => x"ffc348d4",
  1088 => x"99496878",
  1089 => x"c087cd02",
  1090 => x"c702a9ec",
  1091 => x"a9fbc087",
  1092 => x"87cdff05",
  1093 => x"c30266d0",
  1094 => x"7a97c087",
  1095 => x"05a9fbc0",
  1096 => x"4c7387c7",
  1097 => x"c28c0cc0",
  1098 => x"744c7387",
  1099 => x"2687c248",
  1100 => x"264c264d",
  1101 => x"1e4f264b",
  1102 => x"c348d4ff",
  1103 => x"496878ff",
  1104 => x"a9b7f0c0",
  1105 => x"c087ca04",
  1106 => x"01a9b7f9",
  1107 => x"f0c087c3",
  1108 => x"b7c1c189",
  1109 => x"87ca04a9",
  1110 => x"a9b7c6c1",
  1111 => x"c087c301",
  1112 => x"487189f7",
  1113 => x"5e0e4f26",
  1114 => x"0e5d5c5b",
  1115 => x"4c7186f4",
  1116 => x"c04bd4ff",
  1117 => x"ffc37e4d",
  1118 => x"bfd0ff7b",
  1119 => x"c0c0c848",
  1120 => x"58a6c898",
  1121 => x"d0029870",
  1122 => x"bfd0ff87",
  1123 => x"c0c0c848",
  1124 => x"58a6c898",
  1125 => x"f0059870",
  1126 => x"48d0ff87",
  1127 => x"d478e1c0",
  1128 => x"87c2fc7b",
  1129 => x"02994970",
  1130 => x"c387c7c1",
  1131 => x"a6c87bff",
  1132 => x"c8786b48",
  1133 => x"fbc04866",
  1134 => x"87c802a8",
  1135 => x"bfd0fac2",
  1136 => x"87eec002",
  1137 => x"99714dc1",
  1138 => x"87e6c002",
  1139 => x"02a9fbc0",
  1140 => x"d1fb87c3",
  1141 => x"7bffc387",
  1142 => x"c6c1496b",
  1143 => x"87cc05a9",
  1144 => x"7b7bffc3",
  1145 => x"6b48a6c8",
  1146 => x"4d49c078",
  1147 => x"ff059971",
  1148 => x"9d7587da",
  1149 => x"87dec105",
  1150 => x"6b7bffc3",
  1151 => x"7bffc34a",
  1152 => x"6b48a6c4",
  1153 => x"c1486e78",
  1154 => x"58a6c480",
  1155 => x"9749a4c8",
  1156 => x"66c84969",
  1157 => x"87da05a9",
  1158 => x"9749a4c9",
  1159 => x"05aa4969",
  1160 => x"a4ca87d0",
  1161 => x"49699749",
  1162 => x"05a966c4",
  1163 => x"4dc187c4",
  1164 => x"66c887d6",
  1165 => x"a8ecc048",
  1166 => x"c887c902",
  1167 => x"fbc04866",
  1168 => x"87c405a8",
  1169 => x"4dc17ec0",
  1170 => x"c87bffc3",
  1171 => x"786b48a6",
  1172 => x"fe029d75",
  1173 => x"d0ff87e2",
  1174 => x"c0c848bf",
  1175 => x"a6c898c0",
  1176 => x"02987058",
  1177 => x"d0ff87d0",
  1178 => x"c0c848bf",
  1179 => x"a6c898c0",
  1180 => x"05987058",
  1181 => x"d0ff87f0",
  1182 => x"78e0c048",
  1183 => x"8ef4486e",
  1184 => x"0e87ecfa",
  1185 => x"5d5c5b5e",
  1186 => x"c486f40e",
  1187 => x"d0ff59a6",
  1188 => x"c0c0c84c",
  1189 => x"c21e6e4b",
  1190 => x"e949d4fa",
  1191 => x"86c487e7",
  1192 => x"c6029870",
  1193 => x"fac287cb",
  1194 => x"6e4dbfd8",
  1195 => x"87f6fa49",
  1196 => x"7058a6c8",
  1197 => x"4966c41e",
  1198 => x"1e7181c8",
  1199 => x"1ef8d0c1",
  1200 => x"87f8f6fe",
  1201 => x"486c86cc",
  1202 => x"a6cc9873",
  1203 => x"02987058",
  1204 => x"486c87cc",
  1205 => x"a6c49873",
  1206 => x"05987058",
  1207 => x"7cc587f4",
  1208 => x"c148d4ff",
  1209 => x"fac278d5",
  1210 => x"c149bfd0",
  1211 => x"4a66c481",
  1212 => x"32c68ac1",
  1213 => x"b0714872",
  1214 => x"7808d4ff",
  1215 => x"9873486c",
  1216 => x"7058a6c4",
  1217 => x"87cc0298",
  1218 => x"9873486c",
  1219 => x"7058a6c4",
  1220 => x"87f40598",
  1221 => x"d4ff7cc4",
  1222 => x"78ffc348",
  1223 => x"9873486c",
  1224 => x"7058a6c4",
  1225 => x"87cc0298",
  1226 => x"9873486c",
  1227 => x"7058a6c4",
  1228 => x"87f40598",
  1229 => x"d4ff7cc5",
  1230 => x"78d3c148",
  1231 => x"486c78c1",
  1232 => x"a6c49873",
  1233 => x"02987058",
  1234 => x"486c87cc",
  1235 => x"a6c49873",
  1236 => x"05987058",
  1237 => x"7cc487f4",
  1238 => x"c2029d75",
  1239 => x"ecc287d1",
  1240 => x"c21e7ef8",
  1241 => x"eb49d4fa",
  1242 => x"86c487c3",
  1243 => x"c5059870",
  1244 => x"c248c087",
  1245 => x"c0c887fd",
  1246 => x"c404adb7",
  1247 => x"c48d4a87",
  1248 => x"c04a7587",
  1249 => x"73486c4d",
  1250 => x"58a6c898",
  1251 => x"cc029870",
  1252 => x"73486c87",
  1253 => x"58a6c898",
  1254 => x"f4059870",
  1255 => x"ff7ccd87",
  1256 => x"d4c148d4",
  1257 => x"c1497278",
  1258 => x"0299718a",
  1259 => x"976e87d9",
  1260 => x"d4ff48bf",
  1261 => x"486e7808",
  1262 => x"a6c480c1",
  1263 => x"c1497258",
  1264 => x"0599718a",
  1265 => x"6c87e7ff",
  1266 => x"c4987348",
  1267 => x"987058a6",
  1268 => x"6c87cd02",
  1269 => x"c4987348",
  1270 => x"987058a6",
  1271 => x"87f3ff05",
  1272 => x"fac27cc4",
  1273 => x"e1e849d4",
  1274 => x"059d7587",
  1275 => x"6c87effd",
  1276 => x"c4987348",
  1277 => x"987058a6",
  1278 => x"6c87cd02",
  1279 => x"c4987348",
  1280 => x"987058a6",
  1281 => x"87f3ff05",
  1282 => x"d4ff7cc5",
  1283 => x"78d3c148",
  1284 => x"486c78c0",
  1285 => x"a6c49873",
  1286 => x"02987058",
  1287 => x"486c87cd",
  1288 => x"a6c49873",
  1289 => x"05987058",
  1290 => x"c487f3ff",
  1291 => x"c248c17c",
  1292 => x"f448c087",
  1293 => x"87f7f38e",
  1294 => x"6e65704f",
  1295 => x"66206465",
  1296 => x"2c656c69",
  1297 => x"616f6c20",
  1298 => x"676e6964",
  1299 => x"2c732520",
  1300 => x"64692820",
  1301 => x"64252078",
  1302 => x"2e2e2e29",
  1303 => x"6f4c000a",
  1304 => x"6e696461",
  1305 => x"2e2e2e67",
  1306 => x"6c694600",
  1307 => x"73252065",
  1308 => x"2080000a",
  1309 => x"6b636142",
  1310 => x"616f4c00",
  1311 => x"2e2a2064",
  1312 => x"203a0020",
  1313 => x"42208000",
  1314 => x"006b6361",
  1315 => x"78452080",
  1316 => x"49007469",
  1317 => x"6974696e",
  1318 => x"7a696c61",
  1319 => x"20676e69",
  1320 => x"63204453",
  1321 => x"0a647261",
  1322 => x"76614800",
  1323 => x"44532065",
  1324 => x"4f42000a",
  1325 => x"2020544f",
  1326 => x"4f522020",
  1327 => x"5e0e004d",
  1328 => x"0e5d5c5b",
  1329 => x"c04b711e",
  1330 => x"abb74d4c",
  1331 => x"87e9c004",
  1332 => x"1ee6c5c1",
  1333 => x"c4029d75",
  1334 => x"c24ac087",
  1335 => x"724ac187",
  1336 => x"87c6e849",
  1337 => x"58a686c4",
  1338 => x"056e84c1",
  1339 => x"4c7387c2",
  1340 => x"b77385c1",
  1341 => x"d7ff06ac",
  1342 => x"26486e87",
  1343 => x"0e87f0f0",
  1344 => x"5d5c5b5e",
  1345 => x"4c711e0e",
  1346 => x"e4fac249",
  1347 => x"edfe81bf",
  1348 => x"1e4d7087",
  1349 => x"1ee9d1c1",
  1350 => x"87e0edfe",
  1351 => x"9d7586c8",
  1352 => x"87fcc002",
  1353 => x"4bc8f5c2",
  1354 => x"49cb4a75",
  1355 => x"87dbf2fe",
  1356 => x"91de4974",
  1357 => x"48f8fac2",
  1358 => x"a6c48071",
  1359 => x"ded1c158",
  1360 => x"c8496e48",
  1361 => x"41204aa1",
  1362 => x"f905aa71",
  1363 => x"10511087",
  1364 => x"74511051",
  1365 => x"e9c4c149",
  1366 => x"c8f5c287",
  1367 => x"87e3f449",
  1368 => x"49e4f6c1",
  1369 => x"87e5c7c1",
  1370 => x"87c1c8c1",
  1371 => x"87ffee26",
  1372 => x"711e731e",
  1373 => x"fac2494b",
  1374 => x"fd81bfe4",
  1375 => x"4a7087c0",
  1376 => x"87c4029a",
  1377 => x"87dfe349",
  1378 => x"48e4fac2",
  1379 => x"497378c0",
  1380 => x"ee87e9c1",
  1381 => x"731e87dd",
  1382 => x"c44b711e",
  1383 => x"c1024aa3",
  1384 => x"8ac187c8",
  1385 => x"8a87dc02",
  1386 => x"87f1c002",
  1387 => x"c4c1058a",
  1388 => x"e4fac287",
  1389 => x"fcc002bf",
  1390 => x"88c14887",
  1391 => x"58e8fac2",
  1392 => x"c287f2c0",
  1393 => x"49bfe4fa",
  1394 => x"fac289d0",
  1395 => x"b7c059e8",
  1396 => x"e0c003a9",
  1397 => x"e4fac287",
  1398 => x"d878c048",
  1399 => x"e4fac287",
  1400 => x"80c148bf",
  1401 => x"58e8fac2",
  1402 => x"fac287cb",
  1403 => x"d048bfe4",
  1404 => x"e8fac280",
  1405 => x"c3497358",
  1406 => x"87f7ec87",
  1407 => x"5c5b5e0e",
  1408 => x"86f00e5d",
  1409 => x"c259a6d0",
  1410 => x"c04df8ec",
  1411 => x"48a6c44c",
  1412 => x"fac278c0",
  1413 => x"c048bfe4",
  1414 => x"c106a8b7",
  1415 => x"ecc287c1",
  1416 => x"029848f8",
  1417 => x"c187f8c0",
  1418 => x"c81ee6c5",
  1419 => x"87c70266",
  1420 => x"c048a6c4",
  1421 => x"c487c578",
  1422 => x"78c148a6",
  1423 => x"e24966c4",
  1424 => x"86c487e8",
  1425 => x"84c14d70",
  1426 => x"c14866c4",
  1427 => x"58a6c880",
  1428 => x"bfe4fac2",
  1429 => x"c603acb7",
  1430 => x"059d7587",
  1431 => x"c087c8ff",
  1432 => x"029d754c",
  1433 => x"c187e3c3",
  1434 => x"c81ee6c5",
  1435 => x"87c70266",
  1436 => x"c048a6cc",
  1437 => x"cc87c578",
  1438 => x"78c148a6",
  1439 => x"e14966cc",
  1440 => x"86c487e8",
  1441 => x"026e58a6",
  1442 => x"4987ebc2",
  1443 => x"699781cb",
  1444 => x"0299d049",
  1445 => x"c187d9c1",
  1446 => x"744bf0d5",
  1447 => x"c191cc49",
  1448 => x"c881e4f6",
  1449 => x"7a734aa1",
  1450 => x"ffc381c1",
  1451 => x"de497451",
  1452 => x"f8fac291",
  1453 => x"c285714d",
  1454 => x"c17d97c1",
  1455 => x"e0c049a5",
  1456 => x"c8f5c251",
  1457 => x"d202bf97",
  1458 => x"c284c187",
  1459 => x"f5c24ba5",
  1460 => x"49db4ac8",
  1461 => x"87f3ebfe",
  1462 => x"cd87dbc1",
  1463 => x"51c049a5",
  1464 => x"a5c284c1",
  1465 => x"cb4a6e4b",
  1466 => x"deebfe49",
  1467 => x"87c6c187",
  1468 => x"91cc4974",
  1469 => x"81e4f6c1",
  1470 => x"d3c181c8",
  1471 => x"f5c279ff",
  1472 => x"02bf97c8",
  1473 => x"497487d8",
  1474 => x"84c191de",
  1475 => x"4bf8fac2",
  1476 => x"f5c28371",
  1477 => x"49dd4ac8",
  1478 => x"87efeafe",
  1479 => x"4b7487d8",
  1480 => x"fac293de",
  1481 => x"a3cb83f8",
  1482 => x"c151c049",
  1483 => x"4a6e7384",
  1484 => x"eafe49cb",
  1485 => x"66c487d5",
  1486 => x"c880c148",
  1487 => x"b7c758a6",
  1488 => x"c5c003ac",
  1489 => x"fc056e87",
  1490 => x"b7c787dd",
  1491 => x"d3c003ac",
  1492 => x"de497487",
  1493 => x"f8fac291",
  1494 => x"c151c081",
  1495 => x"acb7c784",
  1496 => x"87edff04",
  1497 => x"48f9f7c1",
  1498 => x"f7c150c0",
  1499 => x"50c248f8",
  1500 => x"48c0f8c1",
  1501 => x"78e2dec1",
  1502 => x"48fcf7c1",
  1503 => x"78f2d1c1",
  1504 => x"48ccf8c1",
  1505 => x"78d6d6c1",
  1506 => x"c04966cc",
  1507 => x"f087f3fb",
  1508 => x"87dbe68e",
  1509 => x"c24a711e",
  1510 => x"725ad4fa",
  1511 => x"87dcf949",
  1512 => x"711e4f26",
  1513 => x"91cc494a",
  1514 => x"81e4f6c1",
  1515 => x"481181c1",
  1516 => x"58d0fac2",
  1517 => x"49a2f0c0",
  1518 => x"87dfe8fe",
  1519 => x"ddd549c0",
  1520 => x"0e4f2687",
  1521 => x"5d5c5b5e",
  1522 => x"7186f00e",
  1523 => x"91cc494c",
  1524 => x"81e4f6c1",
  1525 => x"c47ea1c3",
  1526 => x"fac248a6",
  1527 => x"6e78bfc8",
  1528 => x"c44abf97",
  1529 => x"2b724b66",
  1530 => x"124aa1c1",
  1531 => x"58a6cc48",
  1532 => x"83c19b70",
  1533 => x"699781c2",
  1534 => x"04abb749",
  1535 => x"4bc087c2",
  1536 => x"4abf976e",
  1537 => x"724966c8",
  1538 => x"c4b9ff31",
  1539 => x"4d739966",
  1540 => x"b5713572",
  1541 => x"5dccfac2",
  1542 => x"c348d4ff",
  1543 => x"d0ff78ff",
  1544 => x"c0c848bf",
  1545 => x"a6d098c0",
  1546 => x"02987058",
  1547 => x"d0ff87d0",
  1548 => x"c0c848bf",
  1549 => x"a6c498c0",
  1550 => x"05987058",
  1551 => x"d0ff87f0",
  1552 => x"78e1c048",
  1553 => x"de48d4ff",
  1554 => x"7d0d7078",
  1555 => x"c848750d",
  1556 => x"d4ff28b7",
  1557 => x"48757808",
  1558 => x"ff28b7d0",
  1559 => x"757808d4",
  1560 => x"28b7d848",
  1561 => x"7808d4ff",
  1562 => x"48bfd0ff",
  1563 => x"98c0c0c8",
  1564 => x"7058a6c4",
  1565 => x"87d00298",
  1566 => x"48bfd0ff",
  1567 => x"98c0c0c8",
  1568 => x"7058a6c4",
  1569 => x"87f00598",
  1570 => x"c048d0ff",
  1571 => x"1ec778e0",
  1572 => x"f6c11ec0",
  1573 => x"fac21ee4",
  1574 => x"c149bfcc",
  1575 => x"497487e1",
  1576 => x"87def7c0",
  1577 => x"c6e28ee4",
  1578 => x"1e731e87",
  1579 => x"fc494b71",
  1580 => x"497387d1",
  1581 => x"e187ccfc",
  1582 => x"731e87f9",
  1583 => x"c24b711e",
  1584 => x"d5024aa3",
  1585 => x"058ac187",
  1586 => x"fac287db",
  1587 => x"d402bfe0",
  1588 => x"88c14887",
  1589 => x"58e4fac2",
  1590 => x"fac287cb",
  1591 => x"c148bfe0",
  1592 => x"e4fac280",
  1593 => x"c01ec758",
  1594 => x"e4f6c11e",
  1595 => x"ccfac21e",
  1596 => x"87cb49bf",
  1597 => x"f6c04973",
  1598 => x"8ef487c8",
  1599 => x"0e87f4e0",
  1600 => x"5d5c5b5e",
  1601 => x"86d8ff0e",
  1602 => x"c859a6dc",
  1603 => x"78c048a6",
  1604 => x"78c080c4",
  1605 => x"c280c44d",
  1606 => x"78bfe0fa",
  1607 => x"c348d4ff",
  1608 => x"d0ff78ff",
  1609 => x"c0c848bf",
  1610 => x"a6c498c0",
  1611 => x"02987058",
  1612 => x"d0ff87d0",
  1613 => x"c0c848bf",
  1614 => x"a6c498c0",
  1615 => x"05987058",
  1616 => x"d0ff87f0",
  1617 => x"78e1c048",
  1618 => x"d448d4ff",
  1619 => x"d5ddff78",
  1620 => x"48d4ff87",
  1621 => x"d478ffc3",
  1622 => x"d4ff48a6",
  1623 => x"66d478bf",
  1624 => x"a8fbc048",
  1625 => x"87d3c102",
  1626 => x"4a66f8c0",
  1627 => x"7e6a82c4",
  1628 => x"d1c11e72",
  1629 => x"66c448f9",
  1630 => x"4aa1c849",
  1631 => x"aa714120",
  1632 => x"1087f905",
  1633 => x"c04a2651",
  1634 => x"c84966f8",
  1635 => x"d4dec181",
  1636 => x"c7496a79",
  1637 => x"5166d481",
  1638 => x"1ed81ec1",
  1639 => x"81c8496a",
  1640 => x"87d9dcff",
  1641 => x"66d086c8",
  1642 => x"a8b7c048",
  1643 => x"c187c401",
  1644 => x"d087c84d",
  1645 => x"88c14866",
  1646 => x"d458a6d4",
  1647 => x"f4ca0266",
  1648 => x"66c0c187",
  1649 => x"ca03adb7",
  1650 => x"d4ff87eb",
  1651 => x"78ffc348",
  1652 => x"ff48a6d4",
  1653 => x"d478bfd4",
  1654 => x"c6c14866",
  1655 => x"58a6c488",
  1656 => x"c0029870",
  1657 => x"c94887e6",
  1658 => x"58a6c488",
  1659 => x"c4029870",
  1660 => x"c14887d5",
  1661 => x"58a6c488",
  1662 => x"c1029870",
  1663 => x"c44887e3",
  1664 => x"7058a688",
  1665 => x"fec30298",
  1666 => x"87d3c987",
  1667 => x"c10566d8",
  1668 => x"d4ff87c5",
  1669 => x"78ffc348",
  1670 => x"1eca1ec0",
  1671 => x"93cc4b75",
  1672 => x"8366c0c1",
  1673 => x"6c4ca3c4",
  1674 => x"d0daff49",
  1675 => x"de1ec187",
  1676 => x"ff496c1e",
  1677 => x"d087c6da",
  1678 => x"49a3c886",
  1679 => x"79d4dec1",
  1680 => x"adb766d0",
  1681 => x"c187c504",
  1682 => x"87dac885",
  1683 => x"c14866d0",
  1684 => x"58a6d488",
  1685 => x"ff87cfc8",
  1686 => x"d887cbd9",
  1687 => x"c5c858a6",
  1688 => x"d2dbff87",
  1689 => x"58a6cc87",
  1690 => x"a8b766cc",
  1691 => x"cc87c606",
  1692 => x"66c848a6",
  1693 => x"fedaff78",
  1694 => x"a8ecc087",
  1695 => x"87c7c205",
  1696 => x"c10566d8",
  1697 => x"497587f7",
  1698 => x"f8c091cc",
  1699 => x"a1c48166",
  1700 => x"c14c6a4a",
  1701 => x"66c84aa1",
  1702 => x"7997c252",
  1703 => x"dec181c8",
  1704 => x"d4ff79e2",
  1705 => x"78ffc348",
  1706 => x"ff48a6d4",
  1707 => x"d478bfd4",
  1708 => x"e8c00266",
  1709 => x"fbc04887",
  1710 => x"e0c002a8",
  1711 => x"9766d487",
  1712 => x"ff84c17c",
  1713 => x"ffc348d4",
  1714 => x"48a6d478",
  1715 => x"78bfd4ff",
  1716 => x"c80266d4",
  1717 => x"fbc04887",
  1718 => x"e0ff05a8",
  1719 => x"54e0c087",
  1720 => x"c054c1c2",
  1721 => x"66d07c97",
  1722 => x"c504adb7",
  1723 => x"c585c187",
  1724 => x"66d087f4",
  1725 => x"d488c148",
  1726 => x"e9c558a6",
  1727 => x"e5d6ff87",
  1728 => x"58a6d887",
  1729 => x"c887dfc5",
  1730 => x"66d84866",
  1731 => x"c4c505a8",
  1732 => x"48a6dc87",
  1733 => x"d8ff78c0",
  1734 => x"a6d887dd",
  1735 => x"d6d8ff58",
  1736 => x"a6e4c087",
  1737 => x"a8ecc058",
  1738 => x"87cac005",
  1739 => x"48a6e0c0",
  1740 => x"c07866d4",
  1741 => x"d4ff87c6",
  1742 => x"78ffc348",
  1743 => x"91cc4975",
  1744 => x"4866f8c0",
  1745 => x"a6c48071",
  1746 => x"c3496e58",
  1747 => x"5166d481",
  1748 => x"4966e0c0",
  1749 => x"66d481c1",
  1750 => x"7148c189",
  1751 => x"c1497030",
  1752 => x"c14a6e89",
  1753 => x"97097282",
  1754 => x"486e0979",
  1755 => x"fac250c2",
  1756 => x"d449bfc8",
  1757 => x"9729b766",
  1758 => x"71484a6a",
  1759 => x"a6e8c098",
  1760 => x"c4486e58",
  1761 => x"58a6c880",
  1762 => x"4cbf66c4",
  1763 => x"c84866d8",
  1764 => x"c002a866",
  1765 => x"e0c087c9",
  1766 => x"78c048a6",
  1767 => x"c087c6c0",
  1768 => x"c148a6e0",
  1769 => x"66e0c078",
  1770 => x"1ee0c01e",
  1771 => x"d4ff4974",
  1772 => x"86c887cb",
  1773 => x"c058a6d8",
  1774 => x"c106a8b7",
  1775 => x"66d487da",
  1776 => x"bf66c484",
  1777 => x"81e0c049",
  1778 => x"c14b8974",
  1779 => x"714ac2d2",
  1780 => x"87f7d7fe",
  1781 => x"66dc84c2",
  1782 => x"c080c148",
  1783 => x"c058a6e0",
  1784 => x"c14966e4",
  1785 => x"02a97081",
  1786 => x"c087c9c0",
  1787 => x"c048a6e0",
  1788 => x"87c6c078",
  1789 => x"48a6e0c0",
  1790 => x"e0c078c1",
  1791 => x"66c81e66",
  1792 => x"e0c049bf",
  1793 => x"71897481",
  1794 => x"ff49741e",
  1795 => x"c887eed2",
  1796 => x"a8b7c086",
  1797 => x"87fefe01",
  1798 => x"c00266dc",
  1799 => x"496e87d2",
  1800 => x"66dc81c2",
  1801 => x"c8496e51",
  1802 => x"c3dfc181",
  1803 => x"87cdc079",
  1804 => x"81c2496e",
  1805 => x"c8496e51",
  1806 => x"e9e2c181",
  1807 => x"b766d079",
  1808 => x"c5c004ad",
  1809 => x"c085c187",
  1810 => x"66d087dc",
  1811 => x"d488c148",
  1812 => x"d1c058a6",
  1813 => x"cdd1ff87",
  1814 => x"58a6d887",
  1815 => x"ff87c7c0",
  1816 => x"d887c3d1",
  1817 => x"66d458a6",
  1818 => x"87c9c002",
  1819 => x"b766c0c1",
  1820 => x"d5f504ad",
  1821 => x"adb7c787",
  1822 => x"87dcc003",
  1823 => x"91cc4975",
  1824 => x"8166f8c0",
  1825 => x"6a4aa1c4",
  1826 => x"c852c04a",
  1827 => x"c179c081",
  1828 => x"adb7c785",
  1829 => x"87e4ff04",
  1830 => x"c00266d8",
  1831 => x"f8c087eb",
  1832 => x"d4c14966",
  1833 => x"66f8c081",
  1834 => x"82d5c14a",
  1835 => x"51c252c0",
  1836 => x"4966f8c0",
  1837 => x"c181dcc1",
  1838 => x"c079e2de",
  1839 => x"c14966f8",
  1840 => x"d2c181d8",
  1841 => x"d6c079c5",
  1842 => x"66f8c087",
  1843 => x"81d8c149",
  1844 => x"79ccd2c1",
  1845 => x"4966f8c0",
  1846 => x"c281dcc1",
  1847 => x"c179eddd",
  1848 => x"c04afae2",
  1849 => x"c14966f8",
  1850 => x"797281e8",
  1851 => x"48bfd0ff",
  1852 => x"98c0c0c8",
  1853 => x"7058a6c4",
  1854 => x"d1c00298",
  1855 => x"bfd0ff87",
  1856 => x"c0c0c848",
  1857 => x"58a6c498",
  1858 => x"ff059870",
  1859 => x"d0ff87ef",
  1860 => x"78e0c048",
  1861 => x"ff4866cc",
  1862 => x"d0ff8ed8",
  1863 => x"c71e87d1",
  1864 => x"c11ec01e",
  1865 => x"c21ee4f6",
  1866 => x"49bfccfa",
  1867 => x"c187d0ef",
  1868 => x"c049e4f6",
  1869 => x"f487d6e8",
  1870 => x"1e4f268e",
  1871 => x"c287c6ca",
  1872 => x"c048e8fa",
  1873 => x"48d4ff50",
  1874 => x"c178ffc3",
  1875 => x"fe49d3d2",
  1876 => x"fe87d4d1",
  1877 => x"7087d0de",
  1878 => x"87cd0298",
  1879 => x"87d0ebfe",
  1880 => x"c4029870",
  1881 => x"c24ac187",
  1882 => x"724ac087",
  1883 => x"87c8029a",
  1884 => x"49e9d2c1",
  1885 => x"87efd0fe",
  1886 => x"bff8ebc2",
  1887 => x"c2d4ff49",
  1888 => x"e0fac287",
  1889 => x"c278c048",
  1890 => x"c048ccfa",
  1891 => x"cdfe4978",
  1892 => x"87ddc387",
  1893 => x"c087c2c9",
  1894 => x"ff87e1e7",
  1895 => x"4f2687f6",
  1896 => x"000014b2",
  1897 => x"00000002",
  1898 => x"00002eb8",
  1899 => x"000014ff",
  1900 => x"00000002",
  1901 => x"00002ed6",
  1902 => x"000014ff",
  1903 => x"00000002",
  1904 => x"00002ef4",
  1905 => x"000014ff",
  1906 => x"00000002",
  1907 => x"00002f12",
  1908 => x"000014ff",
  1909 => x"00000002",
  1910 => x"00002f30",
  1911 => x"000014ff",
  1912 => x"00000002",
  1913 => x"00002f4e",
  1914 => x"000014ff",
  1915 => x"00000002",
  1916 => x"00002f6c",
  1917 => x"000014ff",
  1918 => x"00000002",
  1919 => x"00000000",
  1920 => x"000017a2",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00001596",
  1924 => x"d5c11e1e",
  1925 => x"58a6c487",
  1926 => x"1e4f2626",
  1927 => x"f0fe4a71",
  1928 => x"cd78c048",
  1929 => x"c10a7a0a",
  1930 => x"fe49f1f8",
  1931 => x"2687f8cd",
  1932 => x"7465534f",
  1933 => x"6e616820",
  1934 => x"72656c64",
  1935 => x"6e49000a",
  1936 => x"746e6920",
  1937 => x"75727265",
  1938 => x"63207470",
  1939 => x"74736e6f",
  1940 => x"74637572",
  1941 => x"000a726f",
  1942 => x"fef8c11e",
  1943 => x"c6cdfe49",
  1944 => x"d0f8c187",
  1945 => x"87f3fe49",
  1946 => x"fe1e4f26",
  1947 => x"2648bff0",
  1948 => x"f0fe1e4f",
  1949 => x"2678c148",
  1950 => x"f0fe1e4f",
  1951 => x"2678c048",
  1952 => x"4a711e4f",
  1953 => x"a2c47ac0",
  1954 => x"c879c049",
  1955 => x"79c049a2",
  1956 => x"c049a2cc",
  1957 => x"0e4f2679",
  1958 => x"0e5c5b5e",
  1959 => x"4c7186f8",
  1960 => x"cc49a4c8",
  1961 => x"486b4ba4",
  1962 => x"a6c480c1",
  1963 => x"c898cf58",
  1964 => x"486958a6",
  1965 => x"05a866c4",
  1966 => x"486b87d4",
  1967 => x"a6c480c1",
  1968 => x"c898cf58",
  1969 => x"486958a6",
  1970 => x"02a866c4",
  1971 => x"e8fe87ec",
  1972 => x"a4d0c187",
  1973 => x"c4486b49",
  1974 => x"58a6c490",
  1975 => x"66d48170",
  1976 => x"c1486b79",
  1977 => x"58a6c880",
  1978 => x"7b7098cf",
  1979 => x"fd87d2c1",
  1980 => x"8ef887ff",
  1981 => x"4d2687c2",
  1982 => x"4b264c26",
  1983 => x"5e0e4f26",
  1984 => x"0e5d5c5b",
  1985 => x"4d7186f8",
  1986 => x"6d4ca5c4",
  1987 => x"05a86c48",
  1988 => x"48ff87c5",
  1989 => x"fd87e5c0",
  1990 => x"a5d087df",
  1991 => x"c4486c4b",
  1992 => x"58a6c490",
  1993 => x"4b6b8370",
  1994 => x"6c9bffc3",
  1995 => x"c880c148",
  1996 => x"98cf58a6",
  1997 => x"f8fc7c70",
  1998 => x"48497387",
  1999 => x"f5fe8ef8",
  2000 => x"1e731e87",
  2001 => x"f0fc86f8",
  2002 => x"4bbfe087",
  2003 => x"c0e0c049",
  2004 => x"e7c00299",
  2005 => x"c34a7387",
  2006 => x"fec29aff",
  2007 => x"c448bfca",
  2008 => x"58a6c490",
  2009 => x"49dafec2",
  2010 => x"79728170",
  2011 => x"bfcafec2",
  2012 => x"c880c148",
  2013 => x"98cf58a6",
  2014 => x"58cefec2",
  2015 => x"c0d04973",
  2016 => x"f2c00299",
  2017 => x"d2fec287",
  2018 => x"fec248bf",
  2019 => x"02a8bfd6",
  2020 => x"c287e4c0",
  2021 => x"48bfd2fe",
  2022 => x"a6c490c4",
  2023 => x"daffc258",
  2024 => x"e0817049",
  2025 => x"c2786948",
  2026 => x"48bfd2fe",
  2027 => x"a6c880c1",
  2028 => x"c298cf58",
  2029 => x"fa58d6fe",
  2030 => x"a6c487f0",
  2031 => x"87f1fa58",
  2032 => x"f5fc8ef8",
  2033 => x"fec21e87",
  2034 => x"f4fa49ca",
  2035 => x"c1fdc187",
  2036 => x"87c7f949",
  2037 => x"2687f5c3",
  2038 => x"1e731e4f",
  2039 => x"49cafec2",
  2040 => x"7087dbfc",
  2041 => x"aab7c04a",
  2042 => x"87ccc204",
  2043 => x"05aaf0c3",
  2044 => x"c2c287c9",
  2045 => x"78c148c4",
  2046 => x"c387edc1",
  2047 => x"c905aae0",
  2048 => x"c8c2c287",
  2049 => x"c178c148",
  2050 => x"c2c287de",
  2051 => x"c602bfc8",
  2052 => x"a2c0c287",
  2053 => x"7287c24b",
  2054 => x"c4c2c24b",
  2055 => x"e0c002bf",
  2056 => x"c4497387",
  2057 => x"c29129b7",
  2058 => x"7381ccc2",
  2059 => x"c29acf4a",
  2060 => x"7248c192",
  2061 => x"ff4a7030",
  2062 => x"694872ba",
  2063 => x"db797098",
  2064 => x"c4497387",
  2065 => x"c29129b7",
  2066 => x"7381ccc2",
  2067 => x"c29acf4a",
  2068 => x"7248c392",
  2069 => x"484a7030",
  2070 => x"7970b069",
  2071 => x"48c8c2c2",
  2072 => x"c2c278c0",
  2073 => x"78c048c4",
  2074 => x"49cafec2",
  2075 => x"7087cffa",
  2076 => x"aab7c04a",
  2077 => x"87f4fd03",
  2078 => x"87c448c0",
  2079 => x"4c264d26",
  2080 => x"4f264b26",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"724ac01e",
  2100 => x"c291c449",
  2101 => x"c081ccc2",
  2102 => x"d082c179",
  2103 => x"ee04aab7",
  2104 => x"0e4f2687",
  2105 => x"5d5c5b5e",
  2106 => x"f64d710e",
  2107 => x"4a7587cb",
  2108 => x"922ab7c4",
  2109 => x"82ccc2c2",
  2110 => x"9ccf4c75",
  2111 => x"496a94c2",
  2112 => x"c32b744b",
  2113 => x"7448c29b",
  2114 => x"ff4c7030",
  2115 => x"714874bc",
  2116 => x"f57a7098",
  2117 => x"487387db",
  2118 => x"1e87e1fd",
  2119 => x"bfd0ff1e",
  2120 => x"c0c0c848",
  2121 => x"58a6c498",
  2122 => x"d0029870",
  2123 => x"bfd0ff87",
  2124 => x"c0c0c848",
  2125 => x"58a6c498",
  2126 => x"f0059870",
  2127 => x"48d0ff87",
  2128 => x"7178e1c4",
  2129 => x"08d4ff48",
  2130 => x"4866c878",
  2131 => x"7808d4ff",
  2132 => x"1e4f2626",
  2133 => x"c84a711e",
  2134 => x"721e4966",
  2135 => x"87fbfe49",
  2136 => x"d0ff86c4",
  2137 => x"c0c848bf",
  2138 => x"a6c498c0",
  2139 => x"02987058",
  2140 => x"d0ff87d0",
  2141 => x"c0c848bf",
  2142 => x"a6c498c0",
  2143 => x"05987058",
  2144 => x"d0ff87f0",
  2145 => x"78e0c048",
  2146 => x"1e4f2626",
  2147 => x"4b711e73",
  2148 => x"731e66c8",
  2149 => x"a2e0c14a",
  2150 => x"87f7fe49",
  2151 => x"2687c426",
  2152 => x"264c264d",
  2153 => x"1e4f264b",
  2154 => x"bfd0ff1e",
  2155 => x"c0c0c848",
  2156 => x"58a6c498",
  2157 => x"d0029870",
  2158 => x"bfd0ff87",
  2159 => x"c0c0c848",
  2160 => x"58a6c498",
  2161 => x"f0059870",
  2162 => x"48d0ff87",
  2163 => x"7178c9c4",
  2164 => x"08d4ff48",
  2165 => x"4f262678",
  2166 => x"4a711e1e",
  2167 => x"87c7ff49",
  2168 => x"48bfd0ff",
  2169 => x"98c0c0c8",
  2170 => x"7058a6c4",
  2171 => x"87d00298",
  2172 => x"48bfd0ff",
  2173 => x"98c0c0c8",
  2174 => x"7058a6c4",
  2175 => x"87f00598",
  2176 => x"c848d0ff",
  2177 => x"4f262678",
  2178 => x"1e1e731e",
  2179 => x"c0c34b71",
  2180 => x"c302bfe6",
  2181 => x"87ccc387",
  2182 => x"48bfd0ff",
  2183 => x"98c0c0c8",
  2184 => x"7058a6c4",
  2185 => x"87d00298",
  2186 => x"48bfd0ff",
  2187 => x"98c0c0c8",
  2188 => x"7058a6c4",
  2189 => x"87f00598",
  2190 => x"c448d0ff",
  2191 => x"487378c9",
  2192 => x"ffb0e0c0",
  2193 => x"c37808d4",
  2194 => x"c048dac0",
  2195 => x"0266cc78",
  2196 => x"ffc387c5",
  2197 => x"c087c249",
  2198 => x"e2c0c349",
  2199 => x"0266d059",
  2200 => x"d5c587c6",
  2201 => x"87c44ad5",
  2202 => x"4affffcf",
  2203 => x"5ae6c0c3",
  2204 => x"48e6c0c3",
  2205 => x"c42678c1",
  2206 => x"264d2687",
  2207 => x"264b264c",
  2208 => x"5b5e0e4f",
  2209 => x"710e5d5c",
  2210 => x"e2c0c34a",
  2211 => x"9a724cbf",
  2212 => x"4987cb02",
  2213 => x"c9c291c8",
  2214 => x"83714bc2",
  2215 => x"cdc287c4",
  2216 => x"4dc04bc2",
  2217 => x"99744913",
  2218 => x"bfdec0c3",
  2219 => x"ffb87148",
  2220 => x"c17808d4",
  2221 => x"c8852cb7",
  2222 => x"e704adb7",
  2223 => x"dac0c387",
  2224 => x"80c848bf",
  2225 => x"58dec0c3",
  2226 => x"1e87eefe",
  2227 => x"4b711e73",
  2228 => x"029a4a13",
  2229 => x"497287cb",
  2230 => x"1387e6fe",
  2231 => x"f5059a4a",
  2232 => x"87d9fe87",
  2233 => x"c0c31e1e",
  2234 => x"c349bfda",
  2235 => x"c148dac0",
  2236 => x"c0c478a1",
  2237 => x"db03a9b7",
  2238 => x"48d4ff87",
  2239 => x"bfdec0c3",
  2240 => x"dac0c378",
  2241 => x"c0c349bf",
  2242 => x"a1c148da",
  2243 => x"b7c0c478",
  2244 => x"87e504a9",
  2245 => x"48bfd0ff",
  2246 => x"98c0c0c8",
  2247 => x"7058a6c4",
  2248 => x"87d00298",
  2249 => x"48bfd0ff",
  2250 => x"98c0c0c8",
  2251 => x"7058a6c4",
  2252 => x"87f00598",
  2253 => x"c848d0ff",
  2254 => x"e6c0c378",
  2255 => x"2678c048",
  2256 => x"00004f26",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"005f5f00",
  2260 => x"03000000",
  2261 => x"03030003",
  2262 => x"7f140000",
  2263 => x"7f7f147f",
  2264 => x"24000014",
  2265 => x"3a6b6b2e",
  2266 => x"6a4c0012",
  2267 => x"566c1836",
  2268 => x"7e300032",
  2269 => x"3a77594f",
  2270 => x"00004068",
  2271 => x"00030704",
  2272 => x"00000000",
  2273 => x"41633e1c",
  2274 => x"00000000",
  2275 => x"1c3e6341",
  2276 => x"2a080000",
  2277 => x"3e1c1c3e",
  2278 => x"0800082a",
  2279 => x"083e3e08",
  2280 => x"00000008",
  2281 => x"0060e080",
  2282 => x"08000000",
  2283 => x"08080808",
  2284 => x"00000008",
  2285 => x"00606000",
  2286 => x"60400000",
  2287 => x"060c1830",
  2288 => x"3e000103",
  2289 => x"7f4d597f",
  2290 => x"0400003e",
  2291 => x"007f7f06",
  2292 => x"42000000",
  2293 => x"4f597163",
  2294 => x"22000046",
  2295 => x"7f494963",
  2296 => x"1c180036",
  2297 => x"7f7f1316",
  2298 => x"27000010",
  2299 => x"7d454567",
  2300 => x"3c000039",
  2301 => x"79494b7e",
  2302 => x"01000030",
  2303 => x"0f797101",
  2304 => x"36000007",
  2305 => x"7f49497f",
  2306 => x"06000036",
  2307 => x"3f69494f",
  2308 => x"0000001e",
  2309 => x"00666600",
  2310 => x"00000000",
  2311 => x"0066e680",
  2312 => x"08000000",
  2313 => x"22141408",
  2314 => x"14000022",
  2315 => x"14141414",
  2316 => x"22000014",
  2317 => x"08141422",
  2318 => x"02000008",
  2319 => x"0f595103",
  2320 => x"7f3e0006",
  2321 => x"1f555d41",
  2322 => x"7e00001e",
  2323 => x"7f09097f",
  2324 => x"7f00007e",
  2325 => x"7f49497f",
  2326 => x"1c000036",
  2327 => x"4141633e",
  2328 => x"7f000041",
  2329 => x"3e63417f",
  2330 => x"7f00001c",
  2331 => x"4149497f",
  2332 => x"7f000041",
  2333 => x"0109097f",
  2334 => x"3e000001",
  2335 => x"7b49417f",
  2336 => x"7f00007a",
  2337 => x"7f08087f",
  2338 => x"0000007f",
  2339 => x"417f7f41",
  2340 => x"20000000",
  2341 => x"7f404060",
  2342 => x"7f7f003f",
  2343 => x"63361c08",
  2344 => x"7f000041",
  2345 => x"4040407f",
  2346 => x"7f7f0040",
  2347 => x"7f060c06",
  2348 => x"7f7f007f",
  2349 => x"7f180c06",
  2350 => x"3e00007f",
  2351 => x"7f41417f",
  2352 => x"7f00003e",
  2353 => x"0f09097f",
  2354 => x"7f3e0006",
  2355 => x"7e7f6141",
  2356 => x"7f000040",
  2357 => x"7f19097f",
  2358 => x"26000066",
  2359 => x"7b594d6f",
  2360 => x"01000032",
  2361 => x"017f7f01",
  2362 => x"3f000001",
  2363 => x"7f40407f",
  2364 => x"0f00003f",
  2365 => x"3f70703f",
  2366 => x"7f7f000f",
  2367 => x"7f301830",
  2368 => x"6341007f",
  2369 => x"361c1c36",
  2370 => x"03014163",
  2371 => x"067c7c06",
  2372 => x"71610103",
  2373 => x"43474d59",
  2374 => x"00000041",
  2375 => x"41417f7f",
  2376 => x"03010000",
  2377 => x"30180c06",
  2378 => x"00004060",
  2379 => x"7f7f4141",
  2380 => x"0c080000",
  2381 => x"0c060306",
  2382 => x"80800008",
  2383 => x"80808080",
  2384 => x"00000080",
  2385 => x"04070300",
  2386 => x"20000000",
  2387 => x"7c545474",
  2388 => x"7f000078",
  2389 => x"7c44447f",
  2390 => x"38000038",
  2391 => x"4444447c",
  2392 => x"38000000",
  2393 => x"7f44447c",
  2394 => x"3800007f",
  2395 => x"5c54547c",
  2396 => x"04000018",
  2397 => x"05057f7e",
  2398 => x"18000000",
  2399 => x"fca4a4bc",
  2400 => x"7f00007c",
  2401 => x"7c04047f",
  2402 => x"00000078",
  2403 => x"407d3d00",
  2404 => x"80000000",
  2405 => x"7dfd8080",
  2406 => x"7f000000",
  2407 => x"6c38107f",
  2408 => x"00000044",
  2409 => x"407f3f00",
  2410 => x"7c7c0000",
  2411 => x"7c0c180c",
  2412 => x"7c000078",
  2413 => x"7c04047c",
  2414 => x"38000078",
  2415 => x"7c44447c",
  2416 => x"fc000038",
  2417 => x"3c2424fc",
  2418 => x"18000018",
  2419 => x"fc24243c",
  2420 => x"7c0000fc",
  2421 => x"0c04047c",
  2422 => x"48000008",
  2423 => x"7454545c",
  2424 => x"04000020",
  2425 => x"44447f3f",
  2426 => x"3c000000",
  2427 => x"7c40407c",
  2428 => x"1c00007c",
  2429 => x"3c60603c",
  2430 => x"7c3c001c",
  2431 => x"7c603060",
  2432 => x"6c44003c",
  2433 => x"6c381038",
  2434 => x"1c000044",
  2435 => x"3c60e0bc",
  2436 => x"4400001c",
  2437 => x"4c5c7464",
  2438 => x"08000044",
  2439 => x"41773e08",
  2440 => x"00000041",
  2441 => x"007f7f00",
  2442 => x"41000000",
  2443 => x"083e7741",
  2444 => x"01020008",
  2445 => x"02020301",
  2446 => x"7f7f0001",
  2447 => x"7f7f7f7f",
  2448 => x"0808007f",
  2449 => x"3e3e1c1c",
  2450 => x"7f7f7f7f",
  2451 => x"1c1c3e3e",
  2452 => x"10000808",
  2453 => x"187c7c18",
  2454 => x"10000010",
  2455 => x"307c7c30",
  2456 => x"30100010",
  2457 => x"1e786060",
  2458 => x"66420006",
  2459 => x"663c183c",
  2460 => x"38780042",
  2461 => x"6cc6c26a",
  2462 => x"00600038",
  2463 => x"00006000",
  2464 => x"5e0e0060",
  2465 => x"0e5d5c5b",
  2466 => x"c34c711e",
  2467 => x"4bbfeec0",
  2468 => x"48f2c0c3",
  2469 => x"1e7478c0",
  2470 => x"1edddcc2",
  2471 => x"87dce7fd",
  2472 => x"6b9786c8",
  2473 => x"c1029949",
  2474 => x"1ec087c6",
  2475 => x"c348a6c4",
  2476 => x"78bff2c0",
  2477 => x"02ac66c4",
  2478 => x"4dc087c4",
  2479 => x"4dc187c2",
  2480 => x"66c81e75",
  2481 => x"87c0ed49",
  2482 => x"e0c086c8",
  2483 => x"87f1ee49",
  2484 => x"6a4aa3c4",
  2485 => x"87f3ef49",
  2486 => x"c387c9f0",
  2487 => x"48bff2c0",
  2488 => x"c0c380c1",
  2489 => x"83cc58f6",
  2490 => x"99496b97",
  2491 => x"87fafe05",
  2492 => x"bff2c0c3",
  2493 => x"adb7c84d",
  2494 => x"c087d903",
  2495 => x"c0c31e1e",
  2496 => x"ec49bff2",
  2497 => x"86c887c2",
  2498 => x"c187d9ef",
  2499 => x"adb7c885",
  2500 => x"87e7ff04",
  2501 => x"264d2626",
  2502 => x"264b264c",
  2503 => x"6769484f",
  2504 => x"67696c68",
  2505 => x"72207468",
  2506 => x"2520776f",
  2507 => x"4d000a64",
  2508 => x"20756e65",
  2509 => x"69736976",
  2510 => x"20656c62",
  2511 => x"000a6425",
  2512 => x"6c6c6143",
  2513 => x"6b636162",
  2514 => x"0a782520",
  2515 => x"4a711e00",
  2516 => x"5af2c0c3",
  2517 => x"bff6c0c3",
  2518 => x"87e6fc49",
  2519 => x"bff2c0c3",
  2520 => x"c389c149",
  2521 => x"7159fac0",
  2522 => x"2687d7fc",
  2523 => x"c0c11e4f",
  2524 => x"87e4e949",
  2525 => x"48e1ebc2",
  2526 => x"4f2678c0",
  2527 => x"5c5b5e0e",
  2528 => x"86f40e5d",
  2529 => x"c048a6c8",
  2530 => x"7ebfec78",
  2531 => x"c0c380fc",
  2532 => x"c378bfee",
  2533 => x"4dbffac0",
  2534 => x"c74cbfe8",
  2535 => x"87c3e549",
  2536 => x"99c24970",
  2537 => x"c287cf05",
  2538 => x"49bfd9eb",
  2539 => x"996eb9ff",
  2540 => x"c00299c1",
  2541 => x"49c787fd",
  2542 => x"7087e8e4",
  2543 => x"87cd0298",
  2544 => x"c787d6e0",
  2545 => x"87dbe449",
  2546 => x"f3059870",
  2547 => x"e1ebc287",
  2548 => x"dcc21ebf",
  2549 => x"e2fd1eef",
  2550 => x"86c887e2",
  2551 => x"bfe1ebc2",
  2552 => x"c2bac14a",
  2553 => x"c15ae5eb",
  2554 => x"e749a2c0",
  2555 => x"a6c887ea",
  2556 => x"c278c148",
  2557 => x"6e48d9eb",
  2558 => x"e1ebc278",
  2559 => x"dac105bf",
  2560 => x"48a6c487",
  2561 => x"78c0c0c8",
  2562 => x"7ee5ebc2",
  2563 => x"49bf976e",
  2564 => x"80c1486e",
  2565 => x"7158a6c4",
  2566 => x"7087c8e3",
  2567 => x"87c30298",
  2568 => x"c4b466c4",
  2569 => x"b7c14866",
  2570 => x"58a6c828",
  2571 => x"ff059870",
  2572 => x"497487da",
  2573 => x"7199ffc3",
  2574 => x"e549c01e",
  2575 => x"497487cd",
  2576 => x"7129b7c8",
  2577 => x"e549c11e",
  2578 => x"86c887c1",
  2579 => x"e249fdc3",
  2580 => x"fac387d1",
  2581 => x"87cbe249",
  2582 => x"7487e9c9",
  2583 => x"99ffc349",
  2584 => x"712cb7c8",
  2585 => x"029c74b4",
  2586 => x"c8ff87df",
  2587 => x"496e7ebf",
  2588 => x"bfddebc2",
  2589 => x"a9c0c289",
  2590 => x"87c4c003",
  2591 => x"87cf4cc0",
  2592 => x"48ddebc2",
  2593 => x"c6c0786e",
  2594 => x"ddebc287",
  2595 => x"7478c048",
  2596 => x"0599c849",
  2597 => x"f5c387ce",
  2598 => x"87c7e149",
  2599 => x"99c24970",
  2600 => x"87eec002",
  2601 => x"bff6c0c3",
  2602 => x"87c9c002",
  2603 => x"c388c148",
  2604 => x"d858fac0",
  2605 => x"f2c0c387",
  2606 => x"91cc49bf",
  2607 => x"c88166c4",
  2608 => x"bf6e7ea1",
  2609 => x"87c5c002",
  2610 => x"7349ff4b",
  2611 => x"48a6c80f",
  2612 => x"497478c1",
  2613 => x"c00599c4",
  2614 => x"f2c387ce",
  2615 => x"87c3e049",
  2616 => x"99c24970",
  2617 => x"87fec002",
  2618 => x"c348a6c8",
  2619 => x"78bff2c0",
  2620 => x"c14966c8",
  2621 => x"f6c0c389",
  2622 => x"b76e7ebf",
  2623 => x"cac006a9",
  2624 => x"80c14887",
  2625 => x"58fac0c3",
  2626 => x"c887d6c0",
  2627 => x"91cc4966",
  2628 => x"c88166c4",
  2629 => x"bf6e7ea1",
  2630 => x"87c5c002",
  2631 => x"7349fe4b",
  2632 => x"48a6c80f",
  2633 => x"fdc378c1",
  2634 => x"f6deff49",
  2635 => x"c2497087",
  2636 => x"eec00299",
  2637 => x"f6c0c387",
  2638 => x"c9c002bf",
  2639 => x"f6c0c387",
  2640 => x"c078c048",
  2641 => x"c0c387d8",
  2642 => x"cc49bff2",
  2643 => x"8166c491",
  2644 => x"6e7ea1c8",
  2645 => x"c5c002bf",
  2646 => x"49fd4b87",
  2647 => x"a6c80f73",
  2648 => x"c378c148",
  2649 => x"ddff49fa",
  2650 => x"497087f9",
  2651 => x"c10299c2",
  2652 => x"a6c887c0",
  2653 => x"f2c0c348",
  2654 => x"66c878bf",
  2655 => x"c488c148",
  2656 => x"c0c358a6",
  2657 => x"6e48bff6",
  2658 => x"c003a8b7",
  2659 => x"c0c387c9",
  2660 => x"786e48f6",
  2661 => x"c887d6c0",
  2662 => x"91cc4966",
  2663 => x"c88166c4",
  2664 => x"bf6e7ea1",
  2665 => x"87c5c002",
  2666 => x"7349fc4b",
  2667 => x"48a6c80f",
  2668 => x"c0c378c1",
  2669 => x"c04bbff6",
  2670 => x"c006abb7",
  2671 => x"8bc187c9",
  2672 => x"01abb7c0",
  2673 => x"7487f7ff",
  2674 => x"99f0c349",
  2675 => x"87cfc005",
  2676 => x"ff49dac1",
  2677 => x"7087ccdc",
  2678 => x"0299c249",
  2679 => x"c387e8c2",
  2680 => x"7ebfeec0",
  2681 => x"bff6c0c3",
  2682 => x"abb7c04b",
  2683 => x"87d0c006",
  2684 => x"80cc486e",
  2685 => x"c158a6c4",
  2686 => x"abb7c08b",
  2687 => x"87f0ff01",
  2688 => x"4abf976e",
  2689 => x"c0028ac1",
  2690 => x"028a87f7",
  2691 => x"8a87d6c0",
  2692 => x"87cac102",
  2693 => x"eec1058a",
  2694 => x"c84a6e87",
  2695 => x"f4496a82",
  2696 => x"e2c187eb",
  2697 => x"c84b6e87",
  2698 => x"c21e6b83",
  2699 => x"fd1ec0dd",
  2700 => x"c887c9d9",
  2701 => x"c34b6b86",
  2702 => x"49bff6c0",
  2703 => x"c6c10f73",
  2704 => x"c8496e87",
  2705 => x"6948c181",
  2706 => x"c3497030",
  2707 => x"48bfeac0",
  2708 => x"c0c3b871",
  2709 => x"a6c858ee",
  2710 => x"c078c148",
  2711 => x"496e87e9",
  2712 => x"486e81c8",
  2713 => x"a6c880cb",
  2714 => x"9766c458",
  2715 => x"a2c14abf",
  2716 => x"4969974b",
  2717 => x"c004abb7",
  2718 => x"4bc087c2",
  2719 => x"970b66c4",
  2720 => x"a6c80b7b",
  2721 => x"7578c148",
  2722 => x"e9c0029d",
  2723 => x"c0026d87",
  2724 => x"496d87e4",
  2725 => x"87cbd9ff",
  2726 => x"99c14970",
  2727 => x"87cbc002",
  2728 => x"c34ba5c4",
  2729 => x"49bff6c0",
  2730 => x"c80f4b6b",
  2731 => x"c5c00285",
  2732 => x"ff056d87",
  2733 => x"66c887dc",
  2734 => x"87c8c002",
  2735 => x"bff6c0c3",
  2736 => x"87feee49",
  2737 => x"ccf18ef4",
  2738 => x"11125887",
  2739 => x"1c1b1d14",
  2740 => x"91595a23",
  2741 => x"ebf2f594",
  2742 => x"000000f4",
  2743 => x"00000000",
  2744 => x"00000000",
  2745 => x"14125800",
  2746 => x"1c1b1d11",
  2747 => x"94595a23",
  2748 => x"ebf2f591",
  2749 => x"000000f4",
  2750 => x"00002afc",
  2751 => x"50505553",
  2752 => x"2054524f",
  2753 => x"0053454e",
  2754 => x"00001e58",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
