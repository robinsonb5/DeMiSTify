///////////////   GLOBAL DEFINES   ////////////////
	
`define GUEST_TOP guest_top	// substitute guest_top (lowercase) by guest's Mist top module name		
`define DEMISTIFY_JOYBITS 8
