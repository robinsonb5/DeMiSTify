
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e0",x"c1",x"c3",x"87"),
    12 => (x"86",x"c0",x"d0",x"4e"),
    13 => (x"49",x"e0",x"c1",x"c3"),
    14 => (x"48",x"ec",x"ec",x"c2"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"ec",x"ec",x"c2",x"87"),
    21 => (x"e8",x"ec",x"c2",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"f3",x"c1",x"87",x"f7"),
    25 => (x"ec",x"c2",x"87",x"f5"),
    26 => (x"ec",x"c2",x"4d",x"ec"),
    27 => (x"ad",x"74",x"4c",x"ec"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"5c",x"5b",x"5e",x"0e"),
    32 => (x"86",x"f0",x"0e",x"5d"),
    33 => (x"a6",x"c4",x"4c",x"c0"),
    34 => (x"c0",x"78",x"c0",x"48"),
    35 => (x"c0",x"4b",x"a6",x"e4"),
    36 => (x"48",x"49",x"66",x"e0"),
    37 => (x"e4",x"c0",x"80",x"c1"),
    38 => (x"48",x"11",x"58",x"a6"),
    39 => (x"70",x"58",x"a6",x"c4"),
    40 => (x"f6",x"c3",x"02",x"98"),
    41 => (x"02",x"66",x"c4",x"87"),
    42 => (x"c4",x"87",x"c6",x"c3"),
    43 => (x"78",x"c0",x"48",x"a6"),
    44 => (x"f0",x"c0",x"4a",x"6e"),
    45 => (x"da",x"c2",x"02",x"8a"),
    46 => (x"8a",x"f3",x"c0",x"87"),
    47 => (x"87",x"db",x"c2",x"02"),
    48 => (x"dc",x"02",x"8a",x"c1"),
    49 => (x"02",x"8a",x"c8",x"87"),
    50 => (x"c4",x"87",x"c8",x"c2"),
    51 => (x"87",x"d1",x"02",x"8a"),
    52 => (x"c1",x"02",x"8a",x"c3"),
    53 => (x"8a",x"c2",x"87",x"eb"),
    54 => (x"c3",x"87",x"c6",x"02"),
    55 => (x"c9",x"c2",x"05",x"8a"),
    56 => (x"73",x"83",x"c4",x"87"),
    57 => (x"69",x"89",x"c4",x"49"),
    58 => (x"c1",x"02",x"6e",x"7e"),
    59 => (x"a6",x"c8",x"87",x"c8"),
    60 => (x"c4",x"78",x"c0",x"48"),
    61 => (x"cc",x"78",x"c0",x"80"),
    62 => (x"4a",x"6e",x"4d",x"66"),
    63 => (x"cf",x"2a",x"b7",x"dc"),
    64 => (x"c4",x"48",x"6e",x"9a"),
    65 => (x"72",x"58",x"a6",x"30"),
    66 => (x"87",x"c5",x"02",x"9a"),
    67 => (x"c1",x"48",x"a6",x"c8"),
    68 => (x"06",x"aa",x"c9",x"78"),
    69 => (x"f7",x"c0",x"87",x"c5"),
    70 => (x"c0",x"87",x"c3",x"82"),
    71 => (x"66",x"c8",x"82",x"f0"),
    72 => (x"72",x"87",x"c7",x"02"),
    73 => (x"87",x"f3",x"c2",x"49"),
    74 => (x"85",x"c1",x"84",x"c1"),
    75 => (x"04",x"ad",x"b7",x"c8"),
    76 => (x"c1",x"87",x"c7",x"ff"),
    77 => (x"f0",x"c0",x"87",x"cf"),
    78 => (x"87",x"df",x"c2",x"49"),
    79 => (x"c4",x"c1",x"84",x"c1"),
    80 => (x"73",x"83",x"c4",x"87"),
    81 => (x"6a",x"8a",x"c4",x"4a"),
    82 => (x"87",x"db",x"c1",x"49"),
    83 => (x"4c",x"a4",x"49",x"70"),
    84 => (x"c4",x"87",x"f2",x"c0"),
    85 => (x"78",x"c1",x"48",x"a6"),
    86 => (x"c4",x"87",x"ea",x"c0"),
    87 => (x"c4",x"4a",x"73",x"83"),
    88 => (x"c1",x"49",x"6a",x"8a"),
    89 => (x"84",x"c1",x"87",x"f5"),
    90 => (x"49",x"6e",x"87",x"db"),
    91 => (x"d4",x"87",x"ec",x"c1"),
    92 => (x"c0",x"48",x"6e",x"87"),
    93 => (x"c7",x"05",x"a8",x"e5"),
    94 => (x"48",x"a6",x"c4",x"87"),
    95 => (x"87",x"c5",x"78",x"c1"),
    96 => (x"d6",x"c1",x"49",x"6e"),
    97 => (x"66",x"e0",x"c0",x"87"),
    98 => (x"80",x"c1",x"48",x"49"),
    99 => (x"58",x"a6",x"e4",x"c0"),
   100 => (x"a6",x"c4",x"48",x"11"),
   101 => (x"05",x"98",x"70",x"58"),
   102 => (x"74",x"87",x"ca",x"fc"),
   103 => (x"26",x"8e",x"f0",x"48"),
   104 => (x"26",x"4c",x"26",x"4d"),
   105 => (x"0e",x"4f",x"26",x"4b"),
   106 => (x"0e",x"5c",x"5b",x"5e"),
   107 => (x"4c",x"c0",x"4b",x"71"),
   108 => (x"02",x"9a",x"4a",x"13"),
   109 => (x"49",x"72",x"87",x"cd"),
   110 => (x"c1",x"87",x"e0",x"c0"),
   111 => (x"9a",x"4a",x"13",x"84"),
   112 => (x"74",x"87",x"f3",x"05"),
   113 => (x"26",x"4c",x"26",x"48"),
   114 => (x"1e",x"4f",x"26",x"4b"),
   115 => (x"73",x"81",x"48",x"73"),
   116 => (x"87",x"c5",x"02",x"a9"),
   117 => (x"f6",x"05",x"53",x"12"),
   118 => (x"1e",x"4f",x"26",x"87"),
   119 => (x"4a",x"c0",x"ff",x"1e"),
   120 => (x"c0",x"c4",x"48",x"6a"),
   121 => (x"58",x"a6",x"c4",x"98"),
   122 => (x"f3",x"02",x"98",x"70"),
   123 => (x"48",x"7a",x"71",x"87"),
   124 => (x"1e",x"4f",x"26",x"26"),
   125 => (x"d4",x"ff",x"1e",x"73"),
   126 => (x"7b",x"ff",x"c3",x"4b"),
   127 => (x"ff",x"c3",x"4a",x"6b"),
   128 => (x"c8",x"49",x"6b",x"7b"),
   129 => (x"c3",x"b1",x"72",x"32"),
   130 => (x"4a",x"6b",x"7b",x"ff"),
   131 => (x"b2",x"71",x"31",x"c8"),
   132 => (x"6b",x"7b",x"ff",x"c3"),
   133 => (x"72",x"32",x"c8",x"49"),
   134 => (x"c4",x"48",x"71",x"b1"),
   135 => (x"26",x"4d",x"26",x"87"),
   136 => (x"26",x"4b",x"26",x"4c"),
   137 => (x"5b",x"5e",x"0e",x"4f"),
   138 => (x"71",x"0e",x"5d",x"5c"),
   139 => (x"4c",x"d4",x"ff",x"4a"),
   140 => (x"ff",x"c3",x"48",x"72"),
   141 => (x"c2",x"7c",x"70",x"98"),
   142 => (x"05",x"bf",x"ec",x"ec"),
   143 => (x"66",x"d0",x"87",x"c8"),
   144 => (x"d4",x"30",x"c9",x"48"),
   145 => (x"66",x"d0",x"58",x"a6"),
   146 => (x"71",x"29",x"d8",x"49"),
   147 => (x"98",x"ff",x"c3",x"48"),
   148 => (x"66",x"d0",x"7c",x"70"),
   149 => (x"71",x"29",x"d0",x"49"),
   150 => (x"98",x"ff",x"c3",x"48"),
   151 => (x"66",x"d0",x"7c",x"70"),
   152 => (x"71",x"29",x"c8",x"49"),
   153 => (x"98",x"ff",x"c3",x"48"),
   154 => (x"66",x"d0",x"7c",x"70"),
   155 => (x"98",x"ff",x"c3",x"48"),
   156 => (x"49",x"72",x"7c",x"70"),
   157 => (x"48",x"71",x"29",x"d0"),
   158 => (x"70",x"98",x"ff",x"c3"),
   159 => (x"c9",x"4b",x"6c",x"7c"),
   160 => (x"c3",x"4d",x"ff",x"f0"),
   161 => (x"d0",x"05",x"ab",x"ff"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"8d",x"c1",x"4b",x"6c"),
   164 => (x"c3",x"87",x"c6",x"02"),
   165 => (x"f0",x"02",x"ab",x"ff"),
   166 => (x"fd",x"48",x"73",x"87"),
   167 => (x"c0",x"1e",x"87",x"ff"),
   168 => (x"48",x"d4",x"ff",x"49"),
   169 => (x"c1",x"78",x"ff",x"c3"),
   170 => (x"b7",x"c8",x"c3",x"81"),
   171 => (x"87",x"f1",x"04",x"a9"),
   172 => (x"73",x"1e",x"4f",x"26"),
   173 => (x"c4",x"87",x"e7",x"1e"),
   174 => (x"c0",x"4b",x"df",x"f8"),
   175 => (x"f0",x"ff",x"c0",x"1e"),
   176 => (x"fd",x"49",x"f7",x"c1"),
   177 => (x"86",x"c4",x"87",x"df"),
   178 => (x"c0",x"05",x"a8",x"c1"),
   179 => (x"d4",x"ff",x"87",x"ea"),
   180 => (x"78",x"ff",x"c3",x"48"),
   181 => (x"c0",x"c0",x"c0",x"c1"),
   182 => (x"c0",x"1e",x"c0",x"c0"),
   183 => (x"e9",x"c1",x"f0",x"e1"),
   184 => (x"87",x"c1",x"fd",x"49"),
   185 => (x"98",x"70",x"86",x"c4"),
   186 => (x"ff",x"87",x"ca",x"05"),
   187 => (x"ff",x"c3",x"48",x"d4"),
   188 => (x"cb",x"48",x"c1",x"78"),
   189 => (x"87",x"e6",x"fe",x"87"),
   190 => (x"fe",x"05",x"8b",x"c1"),
   191 => (x"48",x"c0",x"87",x"fd"),
   192 => (x"1e",x"87",x"de",x"fc"),
   193 => (x"d4",x"ff",x"1e",x"73"),
   194 => (x"78",x"ff",x"c3",x"48"),
   195 => (x"fa",x"49",x"fe",x"cc"),
   196 => (x"4b",x"d3",x"87",x"d5"),
   197 => (x"ff",x"c0",x"1e",x"c0"),
   198 => (x"49",x"c1",x"c1",x"f0"),
   199 => (x"c4",x"87",x"c6",x"fc"),
   200 => (x"05",x"98",x"70",x"86"),
   201 => (x"d4",x"ff",x"87",x"ca"),
   202 => (x"78",x"ff",x"c3",x"48"),
   203 => (x"87",x"cb",x"48",x"c1"),
   204 => (x"c1",x"87",x"eb",x"fd"),
   205 => (x"db",x"ff",x"05",x"8b"),
   206 => (x"fb",x"48",x"c0",x"87"),
   207 => (x"4d",x"43",x"87",x"e3"),
   208 => (x"4d",x"43",x"00",x"44"),
   209 => (x"20",x"38",x"35",x"44"),
   210 => (x"20",x"0a",x"64",x"25"),
   211 => (x"4d",x"43",x"00",x"20"),
   212 => (x"5f",x"38",x"35",x"44"),
   213 => (x"64",x"25",x"20",x"32"),
   214 => (x"00",x"20",x"20",x"0a"),
   215 => (x"35",x"44",x"4d",x"43"),
   216 => (x"64",x"25",x"20",x"38"),
   217 => (x"00",x"20",x"20",x"0a"),
   218 => (x"43",x"48",x"44",x"53"),
   219 => (x"69",x"6e",x"49",x"20"),
   220 => (x"6c",x"61",x"69",x"74"),
   221 => (x"74",x"61",x"7a",x"69"),
   222 => (x"20",x"6e",x"6f",x"69"),
   223 => (x"6f",x"72",x"72",x"65"),
   224 => (x"00",x"0a",x"21",x"72"),
   225 => (x"5f",x"64",x"6d",x"63"),
   226 => (x"38",x"44",x"4d",x"43"),
   227 => (x"73",x"65",x"72",x"20"),
   228 => (x"73",x"6e",x"6f",x"70"),
   229 => (x"25",x"20",x"3a",x"65"),
   230 => (x"49",x"00",x"0a",x"64"),
   231 => (x"00",x"52",x"52",x"45"),
   232 => (x"00",x"49",x"50",x"53"),
   233 => (x"63",x"20",x"44",x"53"),
   234 => (x"20",x"64",x"72",x"61"),
   235 => (x"65",x"7a",x"69",x"73"),
   236 => (x"20",x"73",x"69",x"20"),
   237 => (x"00",x"0a",x"64",x"25"),
   238 => (x"74",x"69",x"72",x"57"),
   239 => (x"61",x"66",x"20",x"65"),
   240 => (x"64",x"65",x"6c",x"69"),
   241 => (x"5f",x"63",x"00",x"0a"),
   242 => (x"65",x"7a",x"69",x"73"),
   243 => (x"6c",x"75",x"6d",x"5f"),
   244 => (x"25",x"20",x"3a",x"74"),
   245 => (x"72",x"20",x"2c",x"64"),
   246 => (x"5f",x"64",x"61",x"65"),
   247 => (x"6c",x"5f",x"6c",x"62"),
   248 => (x"20",x"3a",x"6e",x"65"),
   249 => (x"20",x"2c",x"64",x"25"),
   250 => (x"7a",x"69",x"73",x"63"),
   251 => (x"25",x"20",x"3a",x"65"),
   252 => (x"4d",x"00",x"0a",x"64"),
   253 => (x"20",x"74",x"6c",x"75"),
   254 => (x"00",x"0a",x"64",x"25"),
   255 => (x"62",x"20",x"64",x"25"),
   256 => (x"6b",x"63",x"6f",x"6c"),
   257 => (x"66",x"6f",x"20",x"73"),
   258 => (x"7a",x"69",x"73",x"20"),
   259 => (x"64",x"25",x"20",x"65"),
   260 => (x"64",x"25",x"00",x"0a"),
   261 => (x"6f",x"6c",x"62",x"20"),
   262 => (x"20",x"73",x"6b",x"63"),
   263 => (x"35",x"20",x"66",x"6f"),
   264 => (x"62",x"20",x"32",x"31"),
   265 => (x"73",x"65",x"74",x"79"),
   266 => (x"5e",x"0e",x"00",x"0a"),
   267 => (x"0e",x"5d",x"5c",x"5b"),
   268 => (x"f9",x"4d",x"d4",x"ff"),
   269 => (x"ea",x"c6",x"87",x"e8"),
   270 => (x"f0",x"e1",x"c0",x"1e"),
   271 => (x"f7",x"49",x"c8",x"c1"),
   272 => (x"4b",x"70",x"87",x"e3"),
   273 => (x"1e",x"c4",x"ce",x"1e"),
   274 => (x"cc",x"87",x"f1",x"f0"),
   275 => (x"02",x"ab",x"c1",x"86"),
   276 => (x"ee",x"fa",x"87",x"c8"),
   277 => (x"c2",x"48",x"c0",x"87"),
   278 => (x"d6",x"f6",x"87",x"ca"),
   279 => (x"cf",x"49",x"70",x"87"),
   280 => (x"c6",x"99",x"ff",x"ff"),
   281 => (x"c8",x"02",x"a9",x"ea"),
   282 => (x"87",x"d7",x"fa",x"87"),
   283 => (x"f3",x"c1",x"48",x"c0"),
   284 => (x"7d",x"ff",x"c3",x"87"),
   285 => (x"f8",x"4c",x"f1",x"c0"),
   286 => (x"98",x"70",x"87",x"f8"),
   287 => (x"87",x"cb",x"c1",x"02"),
   288 => (x"ff",x"c0",x"1e",x"c0"),
   289 => (x"49",x"fa",x"c1",x"f0"),
   290 => (x"c4",x"87",x"da",x"f6"),
   291 => (x"9b",x"4b",x"70",x"86"),
   292 => (x"87",x"ed",x"c0",x"05"),
   293 => (x"1e",x"c2",x"cd",x"1e"),
   294 => (x"c3",x"87",x"e1",x"ef"),
   295 => (x"4b",x"6d",x"7d",x"ff"),
   296 => (x"1e",x"ce",x"cd",x"1e"),
   297 => (x"d0",x"87",x"d5",x"ef"),
   298 => (x"7d",x"ff",x"c3",x"86"),
   299 => (x"73",x"7d",x"7d",x"7d"),
   300 => (x"99",x"c0",x"c1",x"49"),
   301 => (x"c1",x"87",x"c5",x"02"),
   302 => (x"87",x"e8",x"c0",x"48"),
   303 => (x"e3",x"c0",x"48",x"c0"),
   304 => (x"cd",x"1e",x"73",x"87"),
   305 => (x"f3",x"ee",x"1e",x"dc"),
   306 => (x"c2",x"86",x"c8",x"87"),
   307 => (x"87",x"cc",x"05",x"ac"),
   308 => (x"ee",x"1e",x"e8",x"cd"),
   309 => (x"86",x"c4",x"87",x"e6"),
   310 => (x"87",x"c8",x"48",x"c0"),
   311 => (x"fe",x"05",x"8c",x"c1"),
   312 => (x"48",x"c0",x"87",x"d5"),
   313 => (x"0e",x"87",x"f6",x"f4"),
   314 => (x"5d",x"5c",x"5b",x"5e"),
   315 => (x"d0",x"ff",x"1e",x"0e"),
   316 => (x"c0",x"c0",x"c8",x"4d"),
   317 => (x"ec",x"ec",x"c2",x"4b"),
   318 => (x"ce",x"78",x"c1",x"48"),
   319 => (x"e6",x"f2",x"49",x"e0"),
   320 => (x"6d",x"4c",x"c7",x"87"),
   321 => (x"c4",x"98",x"73",x"48"),
   322 => (x"98",x"70",x"58",x"a6"),
   323 => (x"6d",x"87",x"cc",x"02"),
   324 => (x"c4",x"98",x"73",x"48"),
   325 => (x"98",x"70",x"58",x"a6"),
   326 => (x"c2",x"87",x"f4",x"05"),
   327 => (x"87",x"fe",x"f5",x"7d"),
   328 => (x"98",x"73",x"48",x"6d"),
   329 => (x"70",x"58",x"a6",x"c4"),
   330 => (x"87",x"cc",x"02",x"98"),
   331 => (x"98",x"73",x"48",x"6d"),
   332 => (x"70",x"58",x"a6",x"c4"),
   333 => (x"87",x"f4",x"05",x"98"),
   334 => (x"1e",x"c0",x"7d",x"c3"),
   335 => (x"c1",x"d0",x"e5",x"c0"),
   336 => (x"e0",x"f3",x"49",x"c0"),
   337 => (x"c1",x"86",x"c4",x"87"),
   338 => (x"87",x"c1",x"05",x"a8"),
   339 => (x"05",x"ac",x"c2",x"4c"),
   340 => (x"db",x"ce",x"87",x"cb"),
   341 => (x"87",x"cf",x"f1",x"49"),
   342 => (x"d8",x"c1",x"48",x"c0"),
   343 => (x"05",x"8c",x"c1",x"87"),
   344 => (x"fb",x"87",x"e0",x"fe"),
   345 => (x"ec",x"c2",x"87",x"c4"),
   346 => (x"98",x"70",x"58",x"f0"),
   347 => (x"c1",x"87",x"cd",x"05"),
   348 => (x"f0",x"ff",x"c0",x"1e"),
   349 => (x"f2",x"49",x"d0",x"c1"),
   350 => (x"86",x"c4",x"87",x"eb"),
   351 => (x"c3",x"48",x"d4",x"ff"),
   352 => (x"e7",x"c5",x"78",x"ff"),
   353 => (x"f4",x"ec",x"c2",x"87"),
   354 => (x"ce",x"1e",x"70",x"58"),
   355 => (x"eb",x"eb",x"1e",x"e4"),
   356 => (x"6d",x"86",x"c8",x"87"),
   357 => (x"c4",x"98",x"73",x"48"),
   358 => (x"98",x"70",x"58",x"a6"),
   359 => (x"6d",x"87",x"cc",x"02"),
   360 => (x"c4",x"98",x"73",x"48"),
   361 => (x"98",x"70",x"58",x"a6"),
   362 => (x"c2",x"87",x"f4",x"05"),
   363 => (x"48",x"d4",x"ff",x"7d"),
   364 => (x"c1",x"78",x"ff",x"c3"),
   365 => (x"e4",x"f1",x"26",x"48"),
   366 => (x"5b",x"5e",x"0e",x"87"),
   367 => (x"1e",x"0e",x"5d",x"5c"),
   368 => (x"4b",x"c0",x"c0",x"c8"),
   369 => (x"ee",x"c5",x"4c",x"c0"),
   370 => (x"c4",x"4a",x"df",x"cd"),
   371 => (x"d4",x"ff",x"5c",x"a6"),
   372 => (x"7c",x"ff",x"c3",x"4c"),
   373 => (x"fe",x"c3",x"48",x"6c"),
   374 => (x"c0",x"c2",x"05",x"a8"),
   375 => (x"05",x"99",x"71",x"87"),
   376 => (x"ff",x"87",x"e2",x"c0"),
   377 => (x"73",x"48",x"bf",x"d0"),
   378 => (x"58",x"a6",x"c4",x"98"),
   379 => (x"ce",x"02",x"98",x"70"),
   380 => (x"bf",x"d0",x"ff",x"87"),
   381 => (x"c4",x"98",x"73",x"48"),
   382 => (x"98",x"70",x"58",x"a6"),
   383 => (x"ff",x"87",x"f2",x"05"),
   384 => (x"d1",x"c4",x"48",x"d0"),
   385 => (x"48",x"66",x"d4",x"78"),
   386 => (x"06",x"a8",x"b7",x"c0"),
   387 => (x"c3",x"87",x"e0",x"c0"),
   388 => (x"4a",x"6c",x"7c",x"ff"),
   389 => (x"c7",x"02",x"99",x"71"),
   390 => (x"97",x"0a",x"71",x"87"),
   391 => (x"81",x"c1",x"0a",x"7a"),
   392 => (x"c1",x"48",x"66",x"d4"),
   393 => (x"58",x"a6",x"d8",x"88"),
   394 => (x"01",x"a8",x"b7",x"c0"),
   395 => (x"c3",x"87",x"e0",x"ff"),
   396 => (x"71",x"7c",x"7c",x"ff"),
   397 => (x"e1",x"c0",x"05",x"99"),
   398 => (x"bf",x"d0",x"ff",x"87"),
   399 => (x"c4",x"98",x"73",x"48"),
   400 => (x"98",x"70",x"58",x"a6"),
   401 => (x"ff",x"87",x"ce",x"02"),
   402 => (x"73",x"48",x"bf",x"d0"),
   403 => (x"58",x"a6",x"c4",x"98"),
   404 => (x"f2",x"05",x"98",x"70"),
   405 => (x"48",x"d0",x"ff",x"87"),
   406 => (x"4a",x"c1",x"78",x"d0"),
   407 => (x"05",x"8a",x"c1",x"7e"),
   408 => (x"6e",x"87",x"ee",x"fd"),
   409 => (x"f4",x"ee",x"26",x"48"),
   410 => (x"5b",x"5e",x"0e",x"87"),
   411 => (x"71",x"1e",x"0e",x"5c"),
   412 => (x"c0",x"c0",x"c8",x"4a"),
   413 => (x"ff",x"4c",x"c0",x"4b"),
   414 => (x"ff",x"c3",x"48",x"d4"),
   415 => (x"bf",x"d0",x"ff",x"78"),
   416 => (x"c4",x"98",x"73",x"48"),
   417 => (x"98",x"70",x"58",x"a6"),
   418 => (x"ff",x"87",x"ce",x"02"),
   419 => (x"73",x"48",x"bf",x"d0"),
   420 => (x"58",x"a6",x"c4",x"98"),
   421 => (x"f2",x"05",x"98",x"70"),
   422 => (x"48",x"d0",x"ff",x"87"),
   423 => (x"ff",x"78",x"c3",x"c4"),
   424 => (x"ff",x"c3",x"48",x"d4"),
   425 => (x"c0",x"1e",x"72",x"78"),
   426 => (x"d1",x"c1",x"f0",x"ff"),
   427 => (x"87",x"f5",x"ed",x"49"),
   428 => (x"98",x"70",x"86",x"c4"),
   429 => (x"87",x"ee",x"c0",x"05"),
   430 => (x"d4",x"1e",x"c0",x"c8"),
   431 => (x"f8",x"fb",x"49",x"66"),
   432 => (x"70",x"86",x"c4",x"87"),
   433 => (x"bf",x"d0",x"ff",x"4c"),
   434 => (x"c4",x"98",x"73",x"48"),
   435 => (x"98",x"70",x"58",x"a6"),
   436 => (x"ff",x"87",x"ce",x"02"),
   437 => (x"73",x"48",x"bf",x"d0"),
   438 => (x"58",x"a6",x"c4",x"98"),
   439 => (x"f2",x"05",x"98",x"70"),
   440 => (x"48",x"d0",x"ff",x"87"),
   441 => (x"48",x"74",x"78",x"c2"),
   442 => (x"87",x"f3",x"ec",x"26"),
   443 => (x"5c",x"5b",x"5e",x"0e"),
   444 => (x"c0",x"1e",x"0e",x"5d"),
   445 => (x"f0",x"ff",x"c0",x"1e"),
   446 => (x"ec",x"49",x"c9",x"c1"),
   447 => (x"1e",x"d2",x"87",x"e7"),
   448 => (x"49",x"fa",x"ec",x"c2"),
   449 => (x"c8",x"87",x"f2",x"fa"),
   450 => (x"c1",x"4d",x"c0",x"86"),
   451 => (x"ad",x"b7",x"d2",x"85"),
   452 => (x"c2",x"87",x"f8",x"04"),
   453 => (x"bf",x"97",x"fa",x"ec"),
   454 => (x"99",x"c0",x"c3",x"49"),
   455 => (x"05",x"a9",x"c0",x"c1"),
   456 => (x"c2",x"87",x"e7",x"c0"),
   457 => (x"bf",x"97",x"c1",x"ed"),
   458 => (x"c2",x"31",x"d0",x"49"),
   459 => (x"bf",x"97",x"c2",x"ed"),
   460 => (x"72",x"32",x"c8",x"4a"),
   461 => (x"c3",x"ed",x"c2",x"b1"),
   462 => (x"b1",x"4a",x"bf",x"97"),
   463 => (x"ff",x"cf",x"4d",x"71"),
   464 => (x"c1",x"9d",x"ff",x"ff"),
   465 => (x"c2",x"35",x"ca",x"85"),
   466 => (x"ed",x"c2",x"87",x"de"),
   467 => (x"4b",x"bf",x"97",x"c3"),
   468 => (x"9b",x"c6",x"33",x"c1"),
   469 => (x"97",x"c4",x"ed",x"c2"),
   470 => (x"b7",x"c7",x"49",x"bf"),
   471 => (x"c2",x"b3",x"71",x"29"),
   472 => (x"bf",x"97",x"ff",x"ec"),
   473 => (x"98",x"cf",x"48",x"49"),
   474 => (x"c2",x"58",x"a6",x"c4"),
   475 => (x"bf",x"97",x"c0",x"ed"),
   476 => (x"ca",x"9c",x"c3",x"4c"),
   477 => (x"c1",x"ed",x"c2",x"34"),
   478 => (x"c2",x"49",x"bf",x"97"),
   479 => (x"c2",x"b4",x"71",x"31"),
   480 => (x"bf",x"97",x"c2",x"ed"),
   481 => (x"99",x"c0",x"c3",x"49"),
   482 => (x"71",x"29",x"b7",x"c6"),
   483 => (x"70",x"1e",x"74",x"b4"),
   484 => (x"cf",x"1e",x"73",x"1e"),
   485 => (x"e3",x"e3",x"1e",x"c6"),
   486 => (x"c1",x"83",x"c2",x"87"),
   487 => (x"70",x"30",x"73",x"48"),
   488 => (x"f3",x"cf",x"1e",x"4b"),
   489 => (x"87",x"d4",x"e3",x"1e"),
   490 => (x"66",x"d8",x"48",x"c1"),
   491 => (x"58",x"a6",x"dc",x"30"),
   492 => (x"4d",x"49",x"a4",x"c1"),
   493 => (x"1e",x"70",x"95",x"73"),
   494 => (x"fc",x"cf",x"1e",x"75"),
   495 => (x"87",x"fc",x"e2",x"1e"),
   496 => (x"6e",x"86",x"e4",x"c0"),
   497 => (x"b7",x"c0",x"c8",x"48"),
   498 => (x"87",x"d2",x"06",x"a8"),
   499 => (x"48",x"6e",x"35",x"c1"),
   500 => (x"c4",x"28",x"b7",x"c1"),
   501 => (x"c0",x"c8",x"58",x"a6"),
   502 => (x"ff",x"01",x"a8",x"b7"),
   503 => (x"1e",x"75",x"87",x"ee"),
   504 => (x"e2",x"1e",x"d2",x"d0"),
   505 => (x"86",x"c8",x"87",x"d6"),
   506 => (x"e8",x"26",x"48",x"75"),
   507 => (x"5e",x"0e",x"87",x"ef"),
   508 => (x"71",x"0e",x"5c",x"5b"),
   509 => (x"d0",x"4c",x"c0",x"4b"),
   510 => (x"b7",x"c0",x"48",x"66"),
   511 => (x"e3",x"c0",x"06",x"a8"),
   512 => (x"cc",x"4a",x"13",x"87"),
   513 => (x"49",x"bf",x"97",x"66"),
   514 => (x"c1",x"48",x"66",x"cc"),
   515 => (x"58",x"a6",x"d0",x"80"),
   516 => (x"02",x"aa",x"b7",x"71"),
   517 => (x"48",x"c1",x"87",x"c4"),
   518 => (x"84",x"c1",x"87",x"cc"),
   519 => (x"ac",x"b7",x"66",x"d0"),
   520 => (x"87",x"dd",x"ff",x"04"),
   521 => (x"87",x"c2",x"48",x"c0"),
   522 => (x"4c",x"26",x"4d",x"26"),
   523 => (x"4f",x"26",x"4b",x"26"),
   524 => (x"5c",x"5b",x"5e",x"0e"),
   525 => (x"f5",x"c2",x"0e",x"5d"),
   526 => (x"78",x"c0",x"48",x"e0"),
   527 => (x"49",x"dd",x"ef",x"c0"),
   528 => (x"c2",x"87",x"e4",x"e5"),
   529 => (x"c0",x"1e",x"d8",x"ed"),
   530 => (x"87",x"dd",x"f8",x"49"),
   531 => (x"98",x"70",x"86",x"c4"),
   532 => (x"c0",x"87",x"cc",x"05"),
   533 => (x"e5",x"49",x"c9",x"ec"),
   534 => (x"48",x"c0",x"87",x"cd"),
   535 => (x"c0",x"87",x"e7",x"ca"),
   536 => (x"e5",x"49",x"ea",x"ef"),
   537 => (x"4b",x"c0",x"87",x"c1"),
   538 => (x"48",x"d8",x"fa",x"c2"),
   539 => (x"1e",x"c8",x"78",x"c1"),
   540 => (x"1e",x"c1",x"f0",x"c0"),
   541 => (x"49",x"ce",x"ee",x"c2"),
   542 => (x"c8",x"87",x"f3",x"fd"),
   543 => (x"05",x"98",x"70",x"86"),
   544 => (x"fa",x"c2",x"87",x"c6"),
   545 => (x"78",x"c0",x"48",x"d8"),
   546 => (x"f0",x"c0",x"1e",x"c8"),
   547 => (x"ee",x"c2",x"1e",x"ca"),
   548 => (x"d9",x"fd",x"49",x"ea"),
   549 => (x"70",x"86",x"c8",x"87"),
   550 => (x"87",x"c6",x"05",x"98"),
   551 => (x"48",x"d8",x"fa",x"c2"),
   552 => (x"fa",x"c2",x"78",x"c0"),
   553 => (x"c0",x"1e",x"bf",x"d8"),
   554 => (x"ff",x"1e",x"d3",x"f0"),
   555 => (x"c8",x"87",x"cd",x"df"),
   556 => (x"d8",x"fa",x"c2",x"86"),
   557 => (x"f7",x"c1",x"02",x"bf"),
   558 => (x"d6",x"f5",x"c2",x"87"),
   559 => (x"1e",x"49",x"bf",x"9f"),
   560 => (x"49",x"d6",x"f5",x"c2"),
   561 => (x"a0",x"c2",x"f8",x"48"),
   562 => (x"d0",x"1e",x"71",x"89"),
   563 => (x"1e",x"c0",x"c8",x"1e"),
   564 => (x"1e",x"fb",x"ec",x"c0"),
   565 => (x"87",x"e4",x"de",x"ff"),
   566 => (x"f4",x"c2",x"86",x"d4"),
   567 => (x"c2",x"4b",x"bf",x"de"),
   568 => (x"bf",x"9f",x"d6",x"f5"),
   569 => (x"ea",x"d6",x"c5",x"4a"),
   570 => (x"c8",x"c0",x"05",x"aa"),
   571 => (x"de",x"f4",x"c2",x"87"),
   572 => (x"d4",x"c0",x"4b",x"bf"),
   573 => (x"d5",x"e9",x"ca",x"87"),
   574 => (x"cc",x"c0",x"02",x"aa"),
   575 => (x"dd",x"ec",x"c0",x"87"),
   576 => (x"87",x"e3",x"e2",x"49"),
   577 => (x"fd",x"c7",x"48",x"c0"),
   578 => (x"c0",x"1e",x"73",x"87"),
   579 => (x"ff",x"1e",x"f8",x"ed"),
   580 => (x"c2",x"87",x"e9",x"dd"),
   581 => (x"73",x"1e",x"d8",x"ed"),
   582 => (x"87",x"cd",x"f5",x"49"),
   583 => (x"98",x"70",x"86",x"cc"),
   584 => (x"87",x"c5",x"c0",x"05"),
   585 => (x"dd",x"c7",x"48",x"c0"),
   586 => (x"d0",x"ee",x"c0",x"87"),
   587 => (x"87",x"f7",x"e1",x"49"),
   588 => (x"1e",x"e6",x"f0",x"c0"),
   589 => (x"87",x"c4",x"dd",x"ff"),
   590 => (x"f0",x"c0",x"1e",x"c8"),
   591 => (x"ee",x"c2",x"1e",x"fe"),
   592 => (x"e9",x"fa",x"49",x"ea"),
   593 => (x"70",x"86",x"cc",x"87"),
   594 => (x"c9",x"c0",x"05",x"98"),
   595 => (x"e0",x"f5",x"c2",x"87"),
   596 => (x"c0",x"78",x"c1",x"48"),
   597 => (x"1e",x"c8",x"87",x"e4"),
   598 => (x"1e",x"c7",x"f1",x"c0"),
   599 => (x"49",x"ce",x"ee",x"c2"),
   600 => (x"c8",x"87",x"cb",x"fa"),
   601 => (x"02",x"98",x"70",x"86"),
   602 => (x"c0",x"87",x"cf",x"c0"),
   603 => (x"ff",x"1e",x"f7",x"ee"),
   604 => (x"c4",x"87",x"c9",x"dc"),
   605 => (x"c6",x"48",x"c0",x"86"),
   606 => (x"f5",x"c2",x"87",x"cc"),
   607 => (x"49",x"bf",x"97",x"d6"),
   608 => (x"05",x"a9",x"d5",x"c1"),
   609 => (x"c2",x"87",x"cd",x"c0"),
   610 => (x"bf",x"97",x"d7",x"f5"),
   611 => (x"a9",x"ea",x"c2",x"49"),
   612 => (x"87",x"c5",x"c0",x"02"),
   613 => (x"ed",x"c5",x"48",x"c0"),
   614 => (x"d8",x"ed",x"c2",x"87"),
   615 => (x"c3",x"4c",x"bf",x"97"),
   616 => (x"c0",x"02",x"ac",x"e9"),
   617 => (x"eb",x"c3",x"87",x"cc"),
   618 => (x"c5",x"c0",x"02",x"ac"),
   619 => (x"c5",x"48",x"c0",x"87"),
   620 => (x"ed",x"c2",x"87",x"d4"),
   621 => (x"49",x"bf",x"97",x"e3"),
   622 => (x"cc",x"c0",x"05",x"99"),
   623 => (x"e4",x"ed",x"c2",x"87"),
   624 => (x"c2",x"49",x"bf",x"97"),
   625 => (x"c5",x"c0",x"02",x"a9"),
   626 => (x"c4",x"48",x"c0",x"87"),
   627 => (x"ed",x"c2",x"87",x"f8"),
   628 => (x"48",x"bf",x"97",x"e5"),
   629 => (x"58",x"dc",x"f5",x"c2"),
   630 => (x"c1",x"4a",x"49",x"70"),
   631 => (x"e0",x"f5",x"c2",x"8a"),
   632 => (x"71",x"1e",x"72",x"5a"),
   633 => (x"d0",x"f1",x"c0",x"1e"),
   634 => (x"cf",x"da",x"ff",x"1e"),
   635 => (x"c2",x"86",x"cc",x"87"),
   636 => (x"bf",x"97",x"e6",x"ed"),
   637 => (x"c2",x"81",x"73",x"49"),
   638 => (x"bf",x"97",x"e7",x"ed"),
   639 => (x"35",x"c8",x"4d",x"4a"),
   640 => (x"f9",x"c2",x"85",x"71"),
   641 => (x"ed",x"c2",x"5d",x"f8"),
   642 => (x"48",x"bf",x"97",x"e8"),
   643 => (x"58",x"cc",x"fa",x"c2"),
   644 => (x"bf",x"e0",x"f5",x"c2"),
   645 => (x"87",x"dc",x"c2",x"02"),
   646 => (x"ef",x"c0",x"1e",x"c8"),
   647 => (x"ee",x"c2",x"1e",x"d4"),
   648 => (x"c9",x"f7",x"49",x"ea"),
   649 => (x"70",x"86",x"c8",x"87"),
   650 => (x"c5",x"c0",x"02",x"98"),
   651 => (x"c3",x"48",x"c0",x"87"),
   652 => (x"f5",x"c2",x"87",x"d4"),
   653 => (x"48",x"4a",x"bf",x"d8"),
   654 => (x"f5",x"c2",x"30",x"c4"),
   655 => (x"fa",x"c2",x"58",x"e8"),
   656 => (x"ed",x"c2",x"5a",x"c8"),
   657 => (x"49",x"bf",x"97",x"fd"),
   658 => (x"ed",x"c2",x"31",x"c8"),
   659 => (x"4b",x"bf",x"97",x"fc"),
   660 => (x"ed",x"c2",x"49",x"a1"),
   661 => (x"4b",x"bf",x"97",x"fe"),
   662 => (x"a1",x"73",x"33",x"d0"),
   663 => (x"ff",x"ed",x"c2",x"49"),
   664 => (x"d8",x"4b",x"bf",x"97"),
   665 => (x"49",x"a1",x"73",x"33"),
   666 => (x"59",x"d0",x"fa",x"c2"),
   667 => (x"bf",x"c8",x"fa",x"c2"),
   668 => (x"f4",x"f9",x"c2",x"91"),
   669 => (x"f9",x"c2",x"81",x"bf"),
   670 => (x"ee",x"c2",x"59",x"fc"),
   671 => (x"4b",x"bf",x"97",x"c5"),
   672 => (x"ee",x"c2",x"33",x"c8"),
   673 => (x"4c",x"bf",x"97",x"c4"),
   674 => (x"ee",x"c2",x"4b",x"a3"),
   675 => (x"4c",x"bf",x"97",x"c6"),
   676 => (x"a3",x"74",x"34",x"d0"),
   677 => (x"c7",x"ee",x"c2",x"4b"),
   678 => (x"cf",x"4c",x"bf",x"97"),
   679 => (x"74",x"34",x"d8",x"9c"),
   680 => (x"fa",x"c2",x"4b",x"a3"),
   681 => (x"8b",x"c2",x"5b",x"c0"),
   682 => (x"fa",x"c2",x"92",x"73"),
   683 => (x"a1",x"72",x"48",x"c0"),
   684 => (x"87",x"cb",x"c1",x"78"),
   685 => (x"97",x"ea",x"ed",x"c2"),
   686 => (x"31",x"c8",x"49",x"bf"),
   687 => (x"97",x"e9",x"ed",x"c2"),
   688 => (x"49",x"a1",x"4a",x"bf"),
   689 => (x"59",x"e8",x"f5",x"c2"),
   690 => (x"ff",x"c7",x"31",x"c5"),
   691 => (x"c2",x"29",x"c9",x"81"),
   692 => (x"c2",x"59",x"c8",x"fa"),
   693 => (x"bf",x"97",x"ef",x"ed"),
   694 => (x"c2",x"32",x"c8",x"4a"),
   695 => (x"bf",x"97",x"ee",x"ed"),
   696 => (x"c2",x"4a",x"a2",x"4b"),
   697 => (x"c2",x"5a",x"d0",x"fa"),
   698 => (x"92",x"bf",x"c8",x"fa"),
   699 => (x"fa",x"c2",x"82",x"75"),
   700 => (x"f9",x"c2",x"5a",x"c4"),
   701 => (x"78",x"c0",x"48",x"fc"),
   702 => (x"48",x"f8",x"f9",x"c2"),
   703 => (x"c0",x"78",x"a1",x"72"),
   704 => (x"87",x"e3",x"cd",x"49"),
   705 => (x"df",x"f4",x"48",x"c1"),
   706 => (x"61",x"65",x"52",x"87"),
   707 => (x"66",x"6f",x"20",x"64"),
   708 => (x"52",x"42",x"4d",x"20"),
   709 => (x"69",x"61",x"66",x"20"),
   710 => (x"0a",x"64",x"65",x"6c"),
   711 => (x"20",x"6f",x"4e",x"00"),
   712 => (x"74",x"72",x"61",x"70"),
   713 => (x"6f",x"69",x"74",x"69"),
   714 => (x"69",x"73",x"20",x"6e"),
   715 => (x"74",x"61",x"6e",x"67"),
   716 => (x"20",x"65",x"72",x"75"),
   717 => (x"6e",x"75",x"6f",x"66"),
   718 => (x"4d",x"00",x"0a",x"64"),
   719 => (x"69",x"73",x"52",x"42"),
   720 => (x"20",x"3a",x"65",x"7a"),
   721 => (x"20",x"2c",x"64",x"25"),
   722 => (x"74",x"72",x"61",x"70"),
   723 => (x"6f",x"69",x"74",x"69"),
   724 => (x"7a",x"69",x"73",x"6e"),
   725 => (x"25",x"20",x"3a",x"65"),
   726 => (x"6f",x"20",x"2c",x"64"),
   727 => (x"65",x"73",x"66",x"66"),
   728 => (x"66",x"6f",x"20",x"74"),
   729 => (x"67",x"69",x"73",x"20"),
   730 => (x"64",x"25",x"20",x"3a"),
   731 => (x"69",x"73",x"20",x"2c"),
   732 => (x"78",x"30",x"20",x"67"),
   733 => (x"00",x"0a",x"78",x"25"),
   734 => (x"64",x"61",x"65",x"52"),
   735 => (x"20",x"67",x"6e",x"69"),
   736 => (x"74",x"6f",x"6f",x"62"),
   737 => (x"63",x"65",x"73",x"20"),
   738 => (x"20",x"72",x"6f",x"74"),
   739 => (x"00",x"0a",x"64",x"25"),
   740 => (x"64",x"61",x"65",x"52"),
   741 => (x"6f",x"6f",x"62",x"20"),
   742 => (x"65",x"73",x"20",x"74"),
   743 => (x"72",x"6f",x"74",x"63"),
   744 => (x"6f",x"72",x"66",x"20"),
   745 => (x"69",x"66",x"20",x"6d"),
   746 => (x"20",x"74",x"73",x"72"),
   747 => (x"74",x"72",x"61",x"70"),
   748 => (x"6f",x"69",x"74",x"69"),
   749 => (x"55",x"00",x"0a",x"6e"),
   750 => (x"70",x"75",x"73",x"6e"),
   751 => (x"74",x"72",x"6f",x"70"),
   752 => (x"70",x"20",x"64",x"65"),
   753 => (x"69",x"74",x"72",x"61"),
   754 => (x"6e",x"6f",x"69",x"74"),
   755 => (x"70",x"79",x"74",x"20"),
   756 => (x"00",x"0d",x"21",x"65"),
   757 => (x"33",x"54",x"41",x"46"),
   758 => (x"20",x"20",x"20",x"32"),
   759 => (x"61",x"65",x"52",x"00"),
   760 => (x"67",x"6e",x"69",x"64"),
   761 => (x"52",x"42",x"4d",x"20"),
   762 => (x"42",x"4d",x"00",x"0a"),
   763 => (x"75",x"73",x"20",x"52"),
   764 => (x"73",x"65",x"63",x"63"),
   765 => (x"6c",x"75",x"66",x"73"),
   766 => (x"72",x"20",x"79",x"6c"),
   767 => (x"0a",x"64",x"61",x"65"),
   768 => (x"54",x"41",x"46",x"00"),
   769 => (x"20",x"20",x"36",x"31"),
   770 => (x"41",x"46",x"00",x"20"),
   771 => (x"20",x"32",x"33",x"54"),
   772 => (x"50",x"00",x"20",x"20"),
   773 => (x"69",x"74",x"72",x"61"),
   774 => (x"6e",x"6f",x"69",x"74"),
   775 => (x"6e",x"75",x"6f",x"63"),
   776 => (x"64",x"25",x"20",x"74"),
   777 => (x"75",x"48",x"00",x"0a"),
   778 => (x"6e",x"69",x"74",x"6e"),
   779 => (x"6f",x"66",x"20",x"67"),
   780 => (x"69",x"66",x"20",x"72"),
   781 => (x"79",x"73",x"65",x"6c"),
   782 => (x"6d",x"65",x"74",x"73"),
   783 => (x"41",x"46",x"00",x"0a"),
   784 => (x"20",x"32",x"33",x"54"),
   785 => (x"46",x"00",x"20",x"20"),
   786 => (x"36",x"31",x"54",x"41"),
   787 => (x"00",x"20",x"20",x"20"),
   788 => (x"73",x"75",x"6c",x"43"),
   789 => (x"20",x"72",x"65",x"74"),
   790 => (x"65",x"7a",x"69",x"73"),
   791 => (x"64",x"25",x"20",x"3a"),
   792 => (x"6c",x"43",x"20",x"2c"),
   793 => (x"65",x"74",x"73",x"75"),
   794 => (x"61",x"6d",x"20",x"72"),
   795 => (x"20",x"2c",x"6b",x"73"),
   796 => (x"00",x"0a",x"64",x"25"),
   797 => (x"6e",x"65",x"70",x"4f"),
   798 => (x"66",x"20",x"64",x"65"),
   799 => (x"2c",x"65",x"6c",x"69"),
   800 => (x"61",x"6f",x"6c",x"20"),
   801 => (x"67",x"6e",x"69",x"64"),
   802 => (x"0a",x"2e",x"2e",x"2e"),
   803 => (x"6e",x"61",x"43",x"00"),
   804 => (x"6f",x"20",x"74",x"27"),
   805 => (x"20",x"6e",x"65",x"70"),
   806 => (x"00",x"0a",x"73",x"25"),
   807 => (x"5c",x"5b",x"5e",x"0e"),
   808 => (x"4a",x"71",x"0e",x"5d"),
   809 => (x"bf",x"e0",x"f5",x"c2"),
   810 => (x"72",x"87",x"cc",x"02"),
   811 => (x"2b",x"b7",x"c7",x"4b"),
   812 => (x"ff",x"c1",x"4d",x"72"),
   813 => (x"72",x"87",x"ca",x"9d"),
   814 => (x"2b",x"b7",x"c8",x"4b"),
   815 => (x"ff",x"c3",x"4d",x"72"),
   816 => (x"d8",x"ed",x"c2",x"9d"),
   817 => (x"f4",x"f9",x"c2",x"1e"),
   818 => (x"81",x"73",x"49",x"bf"),
   819 => (x"87",x"d9",x"e6",x"71"),
   820 => (x"98",x"70",x"86",x"c4"),
   821 => (x"c0",x"87",x"c5",x"05"),
   822 => (x"87",x"e6",x"c0",x"48"),
   823 => (x"bf",x"e0",x"f5",x"c2"),
   824 => (x"75",x"87",x"d2",x"02"),
   825 => (x"c2",x"91",x"c4",x"49"),
   826 => (x"69",x"81",x"d8",x"ed"),
   827 => (x"ff",x"ff",x"cf",x"4c"),
   828 => (x"cb",x"9c",x"ff",x"ff"),
   829 => (x"c2",x"49",x"75",x"87"),
   830 => (x"d8",x"ed",x"c2",x"91"),
   831 => (x"4c",x"69",x"9f",x"81"),
   832 => (x"e3",x"ec",x"48",x"74"),
   833 => (x"5b",x"5e",x"0e",x"87"),
   834 => (x"f4",x"0e",x"5d",x"5c"),
   835 => (x"c0",x"4c",x"71",x"86"),
   836 => (x"d0",x"fa",x"c2",x"4b"),
   837 => (x"a6",x"c4",x"7e",x"bf"),
   838 => (x"d4",x"fa",x"c2",x"48"),
   839 => (x"a6",x"c8",x"78",x"bf"),
   840 => (x"c2",x"78",x"c0",x"48"),
   841 => (x"48",x"bf",x"e4",x"f5"),
   842 => (x"c2",x"06",x"a8",x"c0"),
   843 => (x"66",x"c8",x"87",x"e3"),
   844 => (x"05",x"99",x"cf",x"49"),
   845 => (x"ed",x"c2",x"87",x"d8"),
   846 => (x"66",x"c8",x"1e",x"d8"),
   847 => (x"80",x"c1",x"48",x"49"),
   848 => (x"e4",x"58",x"a6",x"cc"),
   849 => (x"86",x"c4",x"87",x"e3"),
   850 => (x"4b",x"d8",x"ed",x"c2"),
   851 => (x"e0",x"c0",x"87",x"c3"),
   852 => (x"4a",x"6b",x"97",x"83"),
   853 => (x"e7",x"c1",x"02",x"9a"),
   854 => (x"aa",x"e5",x"c3",x"87"),
   855 => (x"87",x"e0",x"c1",x"02"),
   856 => (x"97",x"49",x"a3",x"cb"),
   857 => (x"99",x"d8",x"49",x"69"),
   858 => (x"87",x"d4",x"c1",x"05"),
   859 => (x"d0",x"ff",x"49",x"73"),
   860 => (x"1e",x"cb",x"87",x"f5"),
   861 => (x"1e",x"66",x"e0",x"c0"),
   862 => (x"f1",x"e9",x"49",x"73"),
   863 => (x"70",x"86",x"c8",x"87"),
   864 => (x"fb",x"c0",x"05",x"98"),
   865 => (x"4a",x"a3",x"dc",x"87"),
   866 => (x"6a",x"49",x"a4",x"c4"),
   867 => (x"49",x"a3",x"da",x"79"),
   868 => (x"9f",x"4d",x"a4",x"c8"),
   869 => (x"c2",x"7d",x"48",x"69"),
   870 => (x"02",x"bf",x"e0",x"f5"),
   871 => (x"a3",x"d4",x"87",x"d3"),
   872 => (x"49",x"69",x"9f",x"49"),
   873 => (x"99",x"ff",x"ff",x"c0"),
   874 => (x"30",x"d0",x"48",x"71"),
   875 => (x"c2",x"58",x"a6",x"c4"),
   876 => (x"6e",x"7e",x"c0",x"87"),
   877 => (x"70",x"80",x"6d",x"48"),
   878 => (x"c1",x"7c",x"c0",x"7d"),
   879 => (x"87",x"c5",x"c1",x"48"),
   880 => (x"c1",x"48",x"66",x"c8"),
   881 => (x"58",x"a6",x"cc",x"80"),
   882 => (x"bf",x"e4",x"f5",x"c2"),
   883 => (x"dd",x"fd",x"04",x"a8"),
   884 => (x"e0",x"f5",x"c2",x"87"),
   885 => (x"ea",x"c0",x"02",x"bf"),
   886 => (x"fa",x"49",x"6e",x"87"),
   887 => (x"a6",x"c4",x"87",x"fe"),
   888 => (x"cf",x"49",x"70",x"58"),
   889 => (x"f8",x"ff",x"ff",x"ff"),
   890 => (x"d6",x"02",x"a9",x"99"),
   891 => (x"c2",x"49",x"70",x"87"),
   892 => (x"d8",x"f5",x"c2",x"89"),
   893 => (x"f9",x"c2",x"91",x"bf"),
   894 => (x"71",x"48",x"bf",x"f8"),
   895 => (x"58",x"a6",x"c8",x"80"),
   896 => (x"c0",x"87",x"db",x"fc"),
   897 => (x"e8",x"8e",x"f4",x"48"),
   898 => (x"73",x"1e",x"87",x"de"),
   899 => (x"6a",x"4a",x"71",x"1e"),
   900 => (x"71",x"81",x"c1",x"49"),
   901 => (x"dc",x"f5",x"c2",x"7a"),
   902 => (x"cb",x"05",x"99",x"bf"),
   903 => (x"4b",x"a2",x"c8",x"87"),
   904 => (x"f7",x"f9",x"49",x"6b"),
   905 => (x"7b",x"49",x"70",x"87"),
   906 => (x"ff",x"e7",x"48",x"c1"),
   907 => (x"1e",x"73",x"1e",x"87"),
   908 => (x"f9",x"c2",x"4b",x"71"),
   909 => (x"c8",x"49",x"bf",x"f8"),
   910 => (x"4a",x"6a",x"4a",x"a3"),
   911 => (x"f5",x"c2",x"8a",x"c2"),
   912 => (x"72",x"92",x"bf",x"d8"),
   913 => (x"f5",x"c2",x"49",x"a1"),
   914 => (x"6b",x"4a",x"bf",x"dc"),
   915 => (x"49",x"a1",x"72",x"9a"),
   916 => (x"71",x"1e",x"66",x"c8"),
   917 => (x"c4",x"87",x"d2",x"e0"),
   918 => (x"05",x"98",x"70",x"86"),
   919 => (x"48",x"c0",x"87",x"c4"),
   920 => (x"48",x"c1",x"87",x"c2"),
   921 => (x"0e",x"87",x"c5",x"e7"),
   922 => (x"0e",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"c0",x"4a",x"71"),
   924 => (x"c0",x"02",x"9a",x"72"),
   925 => (x"a2",x"da",x"87",x"e0"),
   926 => (x"4b",x"69",x"9f",x"49"),
   927 => (x"bf",x"e0",x"f5",x"c2"),
   928 => (x"d4",x"87",x"cf",x"02"),
   929 => (x"69",x"9f",x"49",x"a2"),
   930 => (x"ff",x"c0",x"4c",x"49"),
   931 => (x"34",x"d0",x"9c",x"ff"),
   932 => (x"4c",x"c0",x"87",x"c2"),
   933 => (x"9b",x"73",x"b3",x"74"),
   934 => (x"4a",x"87",x"df",x"02"),
   935 => (x"f5",x"c2",x"8a",x"c2"),
   936 => (x"92",x"49",x"bf",x"d8"),
   937 => (x"bf",x"f8",x"f9",x"c2"),
   938 => (x"c2",x"80",x"72",x"48"),
   939 => (x"71",x"58",x"d8",x"fa"),
   940 => (x"c2",x"30",x"c4",x"48"),
   941 => (x"c0",x"58",x"e8",x"f5"),
   942 => (x"f9",x"c2",x"87",x"e9"),
   943 => (x"c2",x"4b",x"bf",x"fc"),
   944 => (x"c2",x"48",x"d4",x"fa"),
   945 => (x"78",x"bf",x"c0",x"fa"),
   946 => (x"bf",x"e0",x"f5",x"c2"),
   947 => (x"c2",x"87",x"c9",x"02"),
   948 => (x"49",x"bf",x"d8",x"f5"),
   949 => (x"87",x"c7",x"31",x"c4"),
   950 => (x"bf",x"c4",x"fa",x"c2"),
   951 => (x"c2",x"31",x"c4",x"49"),
   952 => (x"c2",x"59",x"e8",x"f5"),
   953 => (x"e5",x"5b",x"d4",x"fa"),
   954 => (x"5e",x"0e",x"87",x"c0"),
   955 => (x"0e",x"5d",x"5c",x"5b"),
   956 => (x"4a",x"71",x"86",x"f4"),
   957 => (x"87",x"de",x"02",x"9a"),
   958 => (x"48",x"d4",x"ed",x"c2"),
   959 => (x"ed",x"c2",x"78",x"c0"),
   960 => (x"fa",x"c2",x"48",x"cc"),
   961 => (x"c2",x"78",x"bf",x"d4"),
   962 => (x"c2",x"48",x"d0",x"ed"),
   963 => (x"78",x"bf",x"d0",x"fa"),
   964 => (x"48",x"c2",x"c3",x"c1"),
   965 => (x"f5",x"c2",x"78",x"c0"),
   966 => (x"c2",x"49",x"bf",x"e4"),
   967 => (x"4a",x"bf",x"d4",x"ed"),
   968 => (x"c4",x"03",x"aa",x"71"),
   969 => (x"49",x"72",x"87",x"cc"),
   970 => (x"c0",x"05",x"99",x"cf"),
   971 => (x"ed",x"c2",x"87",x"e1"),
   972 => (x"ed",x"c2",x"1e",x"d8"),
   973 => (x"c2",x"49",x"bf",x"cc"),
   974 => (x"c1",x"48",x"cc",x"ed"),
   975 => (x"ff",x"71",x"78",x"a1"),
   976 => (x"c4",x"87",x"e6",x"dc"),
   977 => (x"fe",x"c2",x"c1",x"86"),
   978 => (x"d8",x"ed",x"c2",x"48"),
   979 => (x"c1",x"87",x"cc",x"78"),
   980 => (x"48",x"bf",x"fe",x"c2"),
   981 => (x"c1",x"80",x"e0",x"c0"),
   982 => (x"c2",x"58",x"c2",x"c3"),
   983 => (x"48",x"bf",x"d4",x"ed"),
   984 => (x"ed",x"c2",x"80",x"c1"),
   985 => (x"be",x"27",x"58",x"d8"),
   986 => (x"bf",x"00",x"00",x"10"),
   987 => (x"9c",x"4c",x"bf",x"97"),
   988 => (x"87",x"ee",x"c2",x"02"),
   989 => (x"02",x"ac",x"e5",x"c3"),
   990 => (x"c1",x"87",x"e7",x"c2"),
   991 => (x"4b",x"bf",x"fe",x"c2"),
   992 => (x"11",x"49",x"a3",x"cb"),
   993 => (x"05",x"ad",x"cf",x"4d"),
   994 => (x"74",x"87",x"d6",x"c1"),
   995 => (x"c1",x"99",x"df",x"49"),
   996 => (x"c2",x"91",x"cd",x"89"),
   997 => (x"c1",x"81",x"e8",x"f5"),
   998 => (x"51",x"12",x"4a",x"a3"),
   999 => (x"12",x"4a",x"a3",x"c3"),
  1000 => (x"4a",x"a3",x"c5",x"51"),
  1001 => (x"a3",x"c7",x"51",x"12"),
  1002 => (x"c9",x"51",x"12",x"4a"),
  1003 => (x"51",x"12",x"4a",x"a3"),
  1004 => (x"12",x"4a",x"a3",x"ce"),
  1005 => (x"4a",x"a3",x"d0",x"51"),
  1006 => (x"a3",x"d2",x"51",x"12"),
  1007 => (x"d4",x"51",x"12",x"4a"),
  1008 => (x"51",x"12",x"4a",x"a3"),
  1009 => (x"12",x"4a",x"a3",x"d6"),
  1010 => (x"4a",x"a3",x"d8",x"51"),
  1011 => (x"a3",x"dc",x"51",x"12"),
  1012 => (x"de",x"51",x"12",x"4a"),
  1013 => (x"51",x"12",x"4a",x"a3"),
  1014 => (x"48",x"c2",x"c3",x"c1"),
  1015 => (x"c1",x"c1",x"78",x"c1"),
  1016 => (x"c8",x"49",x"75",x"87"),
  1017 => (x"f3",x"c0",x"05",x"99"),
  1018 => (x"d0",x"49",x"75",x"87"),
  1019 => (x"87",x"d0",x"05",x"99"),
  1020 => (x"c0",x"02",x"66",x"dc"),
  1021 => (x"49",x"73",x"87",x"ca"),
  1022 => (x"70",x"0f",x"66",x"dc"),
  1023 => (x"87",x"dc",x"02",x"98"),
  1024 => (x"bf",x"c2",x"c3",x"c1"),
  1025 => (x"87",x"c6",x"c0",x"05"),
  1026 => (x"48",x"e8",x"f5",x"c2"),
  1027 => (x"c3",x"c1",x"50",x"c0"),
  1028 => (x"78",x"c0",x"48",x"c2"),
  1029 => (x"bf",x"fe",x"c2",x"c1"),
  1030 => (x"87",x"dc",x"c2",x"48"),
  1031 => (x"48",x"c2",x"c3",x"c1"),
  1032 => (x"f5",x"c2",x"78",x"c0"),
  1033 => (x"c2",x"49",x"bf",x"e4"),
  1034 => (x"4a",x"bf",x"d4",x"ed"),
  1035 => (x"fb",x"04",x"aa",x"71"),
  1036 => (x"fa",x"c2",x"87",x"f4"),
  1037 => (x"c0",x"05",x"bf",x"d4"),
  1038 => (x"f5",x"c2",x"87",x"c8"),
  1039 => (x"c1",x"02",x"bf",x"e0"),
  1040 => (x"ed",x"c2",x"87",x"f4"),
  1041 => (x"f1",x"49",x"bf",x"d0"),
  1042 => (x"ed",x"c2",x"87",x"d2"),
  1043 => (x"7e",x"70",x"58",x"d4"),
  1044 => (x"bf",x"e0",x"f5",x"c2"),
  1045 => (x"87",x"dd",x"c0",x"02"),
  1046 => (x"ff",x"cf",x"49",x"6e"),
  1047 => (x"99",x"f8",x"ff",x"ff"),
  1048 => (x"c8",x"c0",x"02",x"a9"),
  1049 => (x"48",x"a6",x"c4",x"87"),
  1050 => (x"e6",x"c0",x"78",x"c0"),
  1051 => (x"48",x"a6",x"c4",x"87"),
  1052 => (x"de",x"c0",x"78",x"c1"),
  1053 => (x"cf",x"49",x"6e",x"87"),
  1054 => (x"a9",x"99",x"f8",x"ff"),
  1055 => (x"87",x"c8",x"c0",x"02"),
  1056 => (x"c0",x"48",x"a6",x"c8"),
  1057 => (x"87",x"c5",x"c0",x"78"),
  1058 => (x"c1",x"48",x"a6",x"c8"),
  1059 => (x"48",x"a6",x"c4",x"78"),
  1060 => (x"c4",x"78",x"66",x"c8"),
  1061 => (x"dd",x"c0",x"05",x"66"),
  1062 => (x"c2",x"49",x"6e",x"87"),
  1063 => (x"d8",x"f5",x"c2",x"89"),
  1064 => (x"f9",x"c2",x"91",x"bf"),
  1065 => (x"71",x"48",x"bf",x"f8"),
  1066 => (x"d0",x"ed",x"c2",x"80"),
  1067 => (x"d4",x"ed",x"c2",x"58"),
  1068 => (x"f9",x"78",x"c0",x"48"),
  1069 => (x"48",x"c0",x"87",x"e0"),
  1070 => (x"dd",x"ff",x"8e",x"f4"),
  1071 => (x"00",x"00",x"87",x"ea"),
  1072 => (x"00",x"00",x"00",x"00"),
  1073 => (x"ff",x"1e",x"00",x"00"),
  1074 => (x"ff",x"c3",x"48",x"d4"),
  1075 => (x"99",x"49",x"68",x"78"),
  1076 => (x"c0",x"87",x"c6",x"02"),
  1077 => (x"ee",x"05",x"a9",x"fb"),
  1078 => (x"26",x"48",x"71",x"87"),
  1079 => (x"5b",x"5e",x"0e",x"4f"),
  1080 => (x"4a",x"71",x"0e",x"5c"),
  1081 => (x"d4",x"ff",x"4b",x"c0"),
  1082 => (x"78",x"ff",x"c3",x"48"),
  1083 => (x"02",x"99",x"49",x"68"),
  1084 => (x"c0",x"87",x"c1",x"c1"),
  1085 => (x"c0",x"02",x"a9",x"ec"),
  1086 => (x"fb",x"c0",x"87",x"fa"),
  1087 => (x"f3",x"c0",x"02",x"a9"),
  1088 => (x"b7",x"66",x"cc",x"87"),
  1089 => (x"87",x"cc",x"03",x"ab"),
  1090 => (x"c7",x"02",x"66",x"d0"),
  1091 => (x"97",x"09",x"72",x"87"),
  1092 => (x"82",x"c1",x"09",x"79"),
  1093 => (x"c2",x"02",x"99",x"71"),
  1094 => (x"ff",x"83",x"c1",x"87"),
  1095 => (x"ff",x"c3",x"48",x"d4"),
  1096 => (x"99",x"49",x"68",x"78"),
  1097 => (x"c0",x"87",x"cd",x"02"),
  1098 => (x"c7",x"02",x"a9",x"ec"),
  1099 => (x"a9",x"fb",x"c0",x"87"),
  1100 => (x"87",x"cd",x"ff",x"05"),
  1101 => (x"c3",x"02",x"66",x"d0"),
  1102 => (x"7a",x"97",x"c0",x"87"),
  1103 => (x"05",x"a9",x"fb",x"c0"),
  1104 => (x"4c",x"73",x"87",x"c7"),
  1105 => (x"c2",x"8c",x"0c",x"c0"),
  1106 => (x"74",x"4c",x"73",x"87"),
  1107 => (x"26",x"87",x"c2",x"48"),
  1108 => (x"26",x"4c",x"26",x"4d"),
  1109 => (x"1e",x"4f",x"26",x"4b"),
  1110 => (x"c3",x"48",x"d4",x"ff"),
  1111 => (x"49",x"68",x"78",x"ff"),
  1112 => (x"a9",x"b7",x"f0",x"c0"),
  1113 => (x"c0",x"87",x"ca",x"04"),
  1114 => (x"01",x"a9",x"b7",x"f9"),
  1115 => (x"f0",x"c0",x"87",x"c3"),
  1116 => (x"b7",x"c1",x"c1",x"89"),
  1117 => (x"87",x"ca",x"04",x"a9"),
  1118 => (x"a9",x"b7",x"c6",x"c1"),
  1119 => (x"c0",x"87",x"c3",x"01"),
  1120 => (x"48",x"71",x"89",x"f7"),
  1121 => (x"5e",x"0e",x"4f",x"26"),
  1122 => (x"0e",x"5d",x"5c",x"5b"),
  1123 => (x"4c",x"71",x"86",x"f4"),
  1124 => (x"c0",x"4b",x"d4",x"ff"),
  1125 => (x"ff",x"c3",x"7e",x"4d"),
  1126 => (x"bf",x"d0",x"ff",x"7b"),
  1127 => (x"c0",x"c0",x"c8",x"48"),
  1128 => (x"58",x"a6",x"c8",x"98"),
  1129 => (x"d0",x"02",x"98",x"70"),
  1130 => (x"bf",x"d0",x"ff",x"87"),
  1131 => (x"c0",x"c0",x"c8",x"48"),
  1132 => (x"58",x"a6",x"c8",x"98"),
  1133 => (x"f0",x"05",x"98",x"70"),
  1134 => (x"48",x"d0",x"ff",x"87"),
  1135 => (x"d4",x"78",x"e1",x"c0"),
  1136 => (x"87",x"c2",x"fc",x"7b"),
  1137 => (x"02",x"99",x"49",x"70"),
  1138 => (x"c3",x"87",x"c7",x"c1"),
  1139 => (x"a6",x"c8",x"7b",x"ff"),
  1140 => (x"c8",x"78",x"6b",x"48"),
  1141 => (x"fb",x"c0",x"48",x"66"),
  1142 => (x"87",x"c8",x"02",x"a8"),
  1143 => (x"bf",x"f0",x"fa",x"c2"),
  1144 => (x"87",x"ee",x"c0",x"02"),
  1145 => (x"99",x"71",x"4d",x"c1"),
  1146 => (x"87",x"e6",x"c0",x"02"),
  1147 => (x"02",x"a9",x"fb",x"c0"),
  1148 => (x"d1",x"fb",x"87",x"c3"),
  1149 => (x"7b",x"ff",x"c3",x"87"),
  1150 => (x"c6",x"c1",x"49",x"6b"),
  1151 => (x"87",x"cc",x"05",x"a9"),
  1152 => (x"7b",x"7b",x"ff",x"c3"),
  1153 => (x"6b",x"48",x"a6",x"c8"),
  1154 => (x"4d",x"49",x"c0",x"78"),
  1155 => (x"ff",x"05",x"99",x"71"),
  1156 => (x"9d",x"75",x"87",x"da"),
  1157 => (x"87",x"de",x"c1",x"05"),
  1158 => (x"6b",x"7b",x"ff",x"c3"),
  1159 => (x"7b",x"ff",x"c3",x"4a"),
  1160 => (x"6b",x"48",x"a6",x"c4"),
  1161 => (x"c1",x"48",x"6e",x"78"),
  1162 => (x"58",x"a6",x"c4",x"80"),
  1163 => (x"97",x"49",x"a4",x"c8"),
  1164 => (x"66",x"c8",x"49",x"69"),
  1165 => (x"87",x"da",x"05",x"a9"),
  1166 => (x"97",x"49",x"a4",x"c9"),
  1167 => (x"05",x"aa",x"49",x"69"),
  1168 => (x"a4",x"ca",x"87",x"d0"),
  1169 => (x"49",x"69",x"97",x"49"),
  1170 => (x"05",x"a9",x"66",x"c4"),
  1171 => (x"4d",x"c1",x"87",x"c4"),
  1172 => (x"66",x"c8",x"87",x"d6"),
  1173 => (x"a8",x"ec",x"c0",x"48"),
  1174 => (x"c8",x"87",x"c9",x"02"),
  1175 => (x"fb",x"c0",x"48",x"66"),
  1176 => (x"87",x"c4",x"05",x"a8"),
  1177 => (x"4d",x"c1",x"7e",x"c0"),
  1178 => (x"c8",x"7b",x"ff",x"c3"),
  1179 => (x"78",x"6b",x"48",x"a6"),
  1180 => (x"fe",x"02",x"9d",x"75"),
  1181 => (x"d0",x"ff",x"87",x"e2"),
  1182 => (x"c0",x"c8",x"48",x"bf"),
  1183 => (x"a6",x"c8",x"98",x"c0"),
  1184 => (x"02",x"98",x"70",x"58"),
  1185 => (x"d0",x"ff",x"87",x"d0"),
  1186 => (x"c0",x"c8",x"48",x"bf"),
  1187 => (x"a6",x"c8",x"98",x"c0"),
  1188 => (x"05",x"98",x"70",x"58"),
  1189 => (x"d0",x"ff",x"87",x"f0"),
  1190 => (x"78",x"e0",x"c0",x"48"),
  1191 => (x"8e",x"f4",x"48",x"6e"),
  1192 => (x"0e",x"87",x"ec",x"fa"),
  1193 => (x"5d",x"5c",x"5b",x"5e"),
  1194 => (x"c4",x"86",x"f4",x"0e"),
  1195 => (x"d0",x"ff",x"59",x"a6"),
  1196 => (x"c0",x"c0",x"c8",x"4c"),
  1197 => (x"c2",x"1e",x"6e",x"4b"),
  1198 => (x"e9",x"49",x"f4",x"fa"),
  1199 => (x"86",x"c4",x"87",x"c7"),
  1200 => (x"c6",x"02",x"98",x"70"),
  1201 => (x"fa",x"c2",x"87",x"cb"),
  1202 => (x"6e",x"4d",x"bf",x"f8"),
  1203 => (x"87",x"f6",x"fa",x"49"),
  1204 => (x"70",x"58",x"a6",x"c8"),
  1205 => (x"49",x"66",x"c4",x"1e"),
  1206 => (x"1e",x"71",x"81",x"c8"),
  1207 => (x"1e",x"d8",x"d1",x"c1"),
  1208 => (x"87",x"d8",x"f6",x"fe"),
  1209 => (x"48",x"6c",x"86",x"cc"),
  1210 => (x"a6",x"cc",x"98",x"73"),
  1211 => (x"02",x"98",x"70",x"58"),
  1212 => (x"48",x"6c",x"87",x"cc"),
  1213 => (x"a6",x"c4",x"98",x"73"),
  1214 => (x"05",x"98",x"70",x"58"),
  1215 => (x"7c",x"c5",x"87",x"f4"),
  1216 => (x"c1",x"48",x"d4",x"ff"),
  1217 => (x"fa",x"c2",x"78",x"d5"),
  1218 => (x"c1",x"49",x"bf",x"f0"),
  1219 => (x"4a",x"66",x"c4",x"81"),
  1220 => (x"32",x"c6",x"8a",x"c1"),
  1221 => (x"b0",x"71",x"48",x"72"),
  1222 => (x"78",x"08",x"d4",x"ff"),
  1223 => (x"98",x"73",x"48",x"6c"),
  1224 => (x"70",x"58",x"a6",x"c4"),
  1225 => (x"87",x"cc",x"02",x"98"),
  1226 => (x"98",x"73",x"48",x"6c"),
  1227 => (x"70",x"58",x"a6",x"c4"),
  1228 => (x"87",x"f4",x"05",x"98"),
  1229 => (x"d4",x"ff",x"7c",x"c4"),
  1230 => (x"78",x"ff",x"c3",x"48"),
  1231 => (x"98",x"73",x"48",x"6c"),
  1232 => (x"70",x"58",x"a6",x"c4"),
  1233 => (x"87",x"cc",x"02",x"98"),
  1234 => (x"98",x"73",x"48",x"6c"),
  1235 => (x"70",x"58",x"a6",x"c4"),
  1236 => (x"87",x"f4",x"05",x"98"),
  1237 => (x"d4",x"ff",x"7c",x"c5"),
  1238 => (x"78",x"d3",x"c1",x"48"),
  1239 => (x"48",x"6c",x"78",x"c1"),
  1240 => (x"a6",x"c4",x"98",x"73"),
  1241 => (x"02",x"98",x"70",x"58"),
  1242 => (x"48",x"6c",x"87",x"cc"),
  1243 => (x"a6",x"c4",x"98",x"73"),
  1244 => (x"05",x"98",x"70",x"58"),
  1245 => (x"7c",x"c4",x"87",x"f4"),
  1246 => (x"c2",x"02",x"9d",x"75"),
  1247 => (x"ed",x"c2",x"87",x"d1"),
  1248 => (x"c2",x"1e",x"7e",x"d8"),
  1249 => (x"ea",x"49",x"f4",x"fa"),
  1250 => (x"86",x"c4",x"87",x"e3"),
  1251 => (x"c5",x"05",x"98",x"70"),
  1252 => (x"c2",x"48",x"c0",x"87"),
  1253 => (x"c0",x"c8",x"87",x"fd"),
  1254 => (x"c4",x"04",x"ad",x"b7"),
  1255 => (x"c4",x"8d",x"4a",x"87"),
  1256 => (x"c0",x"4a",x"75",x"87"),
  1257 => (x"73",x"48",x"6c",x"4d"),
  1258 => (x"58",x"a6",x"c8",x"98"),
  1259 => (x"cc",x"02",x"98",x"70"),
  1260 => (x"73",x"48",x"6c",x"87"),
  1261 => (x"58",x"a6",x"c8",x"98"),
  1262 => (x"f4",x"05",x"98",x"70"),
  1263 => (x"ff",x"7c",x"cd",x"87"),
  1264 => (x"d4",x"c1",x"48",x"d4"),
  1265 => (x"c1",x"49",x"72",x"78"),
  1266 => (x"02",x"99",x"71",x"8a"),
  1267 => (x"97",x"6e",x"87",x"d9"),
  1268 => (x"d4",x"ff",x"48",x"bf"),
  1269 => (x"48",x"6e",x"78",x"08"),
  1270 => (x"a6",x"c4",x"80",x"c1"),
  1271 => (x"c1",x"49",x"72",x"58"),
  1272 => (x"05",x"99",x"71",x"8a"),
  1273 => (x"6c",x"87",x"e7",x"ff"),
  1274 => (x"c4",x"98",x"73",x"48"),
  1275 => (x"98",x"70",x"58",x"a6"),
  1276 => (x"6c",x"87",x"cd",x"02"),
  1277 => (x"c4",x"98",x"73",x"48"),
  1278 => (x"98",x"70",x"58",x"a6"),
  1279 => (x"87",x"f3",x"ff",x"05"),
  1280 => (x"fa",x"c2",x"7c",x"c4"),
  1281 => (x"c1",x"e8",x"49",x"f4"),
  1282 => (x"05",x"9d",x"75",x"87"),
  1283 => (x"6c",x"87",x"ef",x"fd"),
  1284 => (x"c4",x"98",x"73",x"48"),
  1285 => (x"98",x"70",x"58",x"a6"),
  1286 => (x"6c",x"87",x"cd",x"02"),
  1287 => (x"c4",x"98",x"73",x"48"),
  1288 => (x"98",x"70",x"58",x"a6"),
  1289 => (x"87",x"f3",x"ff",x"05"),
  1290 => (x"d4",x"ff",x"7c",x"c5"),
  1291 => (x"78",x"d3",x"c1",x"48"),
  1292 => (x"48",x"6c",x"78",x"c0"),
  1293 => (x"a6",x"c4",x"98",x"73"),
  1294 => (x"02",x"98",x"70",x"58"),
  1295 => (x"48",x"6c",x"87",x"cd"),
  1296 => (x"a6",x"c4",x"98",x"73"),
  1297 => (x"05",x"98",x"70",x"58"),
  1298 => (x"c4",x"87",x"f3",x"ff"),
  1299 => (x"c2",x"48",x"c1",x"7c"),
  1300 => (x"f4",x"48",x"c0",x"87"),
  1301 => (x"87",x"f7",x"f3",x"8e"),
  1302 => (x"6e",x"65",x"70",x"4f"),
  1303 => (x"66",x"20",x"64",x"65"),
  1304 => (x"2c",x"65",x"6c",x"69"),
  1305 => (x"61",x"6f",x"6c",x"20"),
  1306 => (x"67",x"6e",x"69",x"64"),
  1307 => (x"2c",x"73",x"25",x"20"),
  1308 => (x"64",x"69",x"28",x"20"),
  1309 => (x"64",x"25",x"20",x"78"),
  1310 => (x"2e",x"2e",x"2e",x"29"),
  1311 => (x"6f",x"4c",x"00",x"0a"),
  1312 => (x"6e",x"69",x"64",x"61"),
  1313 => (x"2e",x"2e",x"2e",x"67"),
  1314 => (x"6c",x"69",x"46",x"00"),
  1315 => (x"73",x"25",x"20",x"65"),
  1316 => (x"20",x"80",x"00",x"0a"),
  1317 => (x"6b",x"63",x"61",x"42"),
  1318 => (x"61",x"6f",x"4c",x"00"),
  1319 => (x"2e",x"2a",x"20",x"64"),
  1320 => (x"20",x"3a",x"00",x"20"),
  1321 => (x"42",x"20",x"80",x"00"),
  1322 => (x"00",x"6b",x"63",x"61"),
  1323 => (x"78",x"45",x"20",x"80"),
  1324 => (x"49",x"00",x"74",x"69"),
  1325 => (x"69",x"74",x"69",x"6e"),
  1326 => (x"7a",x"69",x"6c",x"61"),
  1327 => (x"20",x"67",x"6e",x"69"),
  1328 => (x"63",x"20",x"44",x"53"),
  1329 => (x"0a",x"64",x"72",x"61"),
  1330 => (x"76",x"61",x"48",x"00"),
  1331 => (x"44",x"53",x"20",x"65"),
  1332 => (x"4f",x"42",x"00",x"0a"),
  1333 => (x"20",x"20",x"54",x"4f"),
  1334 => (x"4f",x"52",x"20",x"20"),
  1335 => (x"5e",x"0e",x"00",x"4d"),
  1336 => (x"0e",x"5d",x"5c",x"5b"),
  1337 => (x"c0",x"4b",x"71",x"1e"),
  1338 => (x"ab",x"b7",x"4d",x"4c"),
  1339 => (x"87",x"e9",x"c0",x"04"),
  1340 => (x"1e",x"c6",x"c6",x"c1"),
  1341 => (x"c4",x"02",x"9d",x"75"),
  1342 => (x"c2",x"4a",x"c0",x"87"),
  1343 => (x"72",x"4a",x"c1",x"87"),
  1344 => (x"87",x"e6",x"e7",x"49"),
  1345 => (x"58",x"a6",x"86",x"c4"),
  1346 => (x"05",x"6e",x"84",x"c1"),
  1347 => (x"4c",x"73",x"87",x"c2"),
  1348 => (x"b7",x"73",x"85",x"c1"),
  1349 => (x"d7",x"ff",x"06",x"ac"),
  1350 => (x"26",x"48",x"6e",x"87"),
  1351 => (x"0e",x"87",x"f0",x"f0"),
  1352 => (x"5d",x"5c",x"5b",x"5e"),
  1353 => (x"4c",x"71",x"1e",x"0e"),
  1354 => (x"c4",x"fb",x"c2",x"49"),
  1355 => (x"ed",x"fe",x"81",x"bf"),
  1356 => (x"1e",x"4d",x"70",x"87"),
  1357 => (x"1e",x"c9",x"d2",x"c1"),
  1358 => (x"87",x"c0",x"ed",x"fe"),
  1359 => (x"9d",x"75",x"86",x"c8"),
  1360 => (x"87",x"fc",x"c0",x"02"),
  1361 => (x"4b",x"e8",x"f5",x"c2"),
  1362 => (x"49",x"cb",x"4a",x"75"),
  1363 => (x"87",x"fb",x"f1",x"fe"),
  1364 => (x"91",x"de",x"49",x"74"),
  1365 => (x"48",x"d8",x"fb",x"c2"),
  1366 => (x"a6",x"c4",x"80",x"71"),
  1367 => (x"fe",x"d1",x"c1",x"58"),
  1368 => (x"c8",x"49",x"6e",x"48"),
  1369 => (x"41",x"20",x"4a",x"a1"),
  1370 => (x"f9",x"05",x"aa",x"71"),
  1371 => (x"10",x"51",x"10",x"87"),
  1372 => (x"74",x"51",x"10",x"51"),
  1373 => (x"e9",x"c4",x"c1",x"49"),
  1374 => (x"e8",x"f5",x"c2",x"87"),
  1375 => (x"87",x"e3",x"f4",x"49"),
  1376 => (x"49",x"c4",x"f7",x"c1"),
  1377 => (x"87",x"e5",x"c7",x"c1"),
  1378 => (x"87",x"c1",x"c8",x"c1"),
  1379 => (x"87",x"ff",x"ee",x"26"),
  1380 => (x"71",x"1e",x"73",x"1e"),
  1381 => (x"fb",x"c2",x"49",x"4b"),
  1382 => (x"fd",x"81",x"bf",x"c4"),
  1383 => (x"4a",x"70",x"87",x"c0"),
  1384 => (x"87",x"c4",x"02",x"9a"),
  1385 => (x"87",x"ff",x"e2",x"49"),
  1386 => (x"48",x"c4",x"fb",x"c2"),
  1387 => (x"49",x"73",x"78",x"c0"),
  1388 => (x"ee",x"87",x"e9",x"c1"),
  1389 => (x"73",x"1e",x"87",x"dd"),
  1390 => (x"c4",x"4b",x"71",x"1e"),
  1391 => (x"c1",x"02",x"4a",x"a3"),
  1392 => (x"8a",x"c1",x"87",x"c8"),
  1393 => (x"8a",x"87",x"dc",x"02"),
  1394 => (x"87",x"f1",x"c0",x"02"),
  1395 => (x"c4",x"c1",x"05",x"8a"),
  1396 => (x"c4",x"fb",x"c2",x"87"),
  1397 => (x"fc",x"c0",x"02",x"bf"),
  1398 => (x"88",x"c1",x"48",x"87"),
  1399 => (x"58",x"c8",x"fb",x"c2"),
  1400 => (x"c2",x"87",x"f2",x"c0"),
  1401 => (x"49",x"bf",x"c4",x"fb"),
  1402 => (x"fb",x"c2",x"89",x"d0"),
  1403 => (x"b7",x"c0",x"59",x"c8"),
  1404 => (x"e0",x"c0",x"03",x"a9"),
  1405 => (x"c4",x"fb",x"c2",x"87"),
  1406 => (x"d8",x"78",x"c0",x"48"),
  1407 => (x"c4",x"fb",x"c2",x"87"),
  1408 => (x"80",x"c1",x"48",x"bf"),
  1409 => (x"58",x"c8",x"fb",x"c2"),
  1410 => (x"fb",x"c2",x"87",x"cb"),
  1411 => (x"d0",x"48",x"bf",x"c4"),
  1412 => (x"c8",x"fb",x"c2",x"80"),
  1413 => (x"c3",x"49",x"73",x"58"),
  1414 => (x"87",x"f7",x"ec",x"87"),
  1415 => (x"5c",x"5b",x"5e",x"0e"),
  1416 => (x"86",x"f0",x"0e",x"5d"),
  1417 => (x"c2",x"59",x"a6",x"d0"),
  1418 => (x"c0",x"4d",x"d8",x"ed"),
  1419 => (x"48",x"a6",x"c4",x"4c"),
  1420 => (x"fb",x"c2",x"78",x"c0"),
  1421 => (x"c0",x"48",x"bf",x"c4"),
  1422 => (x"c1",x"06",x"a8",x"b7"),
  1423 => (x"ed",x"c2",x"87",x"c1"),
  1424 => (x"02",x"98",x"48",x"d8"),
  1425 => (x"c1",x"87",x"f8",x"c0"),
  1426 => (x"c8",x"1e",x"c6",x"c6"),
  1427 => (x"87",x"c7",x"02",x"66"),
  1428 => (x"c0",x"48",x"a6",x"c4"),
  1429 => (x"c4",x"87",x"c5",x"78"),
  1430 => (x"78",x"c1",x"48",x"a6"),
  1431 => (x"e2",x"49",x"66",x"c4"),
  1432 => (x"86",x"c4",x"87",x"c8"),
  1433 => (x"84",x"c1",x"4d",x"70"),
  1434 => (x"c1",x"48",x"66",x"c4"),
  1435 => (x"58",x"a6",x"c8",x"80"),
  1436 => (x"bf",x"c4",x"fb",x"c2"),
  1437 => (x"c6",x"03",x"ac",x"b7"),
  1438 => (x"05",x"9d",x"75",x"87"),
  1439 => (x"c0",x"87",x"c8",x"ff"),
  1440 => (x"02",x"9d",x"75",x"4c"),
  1441 => (x"c1",x"87",x"e3",x"c3"),
  1442 => (x"c8",x"1e",x"c6",x"c6"),
  1443 => (x"87",x"c7",x"02",x"66"),
  1444 => (x"c0",x"48",x"a6",x"cc"),
  1445 => (x"cc",x"87",x"c5",x"78"),
  1446 => (x"78",x"c1",x"48",x"a6"),
  1447 => (x"e1",x"49",x"66",x"cc"),
  1448 => (x"86",x"c4",x"87",x"c8"),
  1449 => (x"02",x"6e",x"58",x"a6"),
  1450 => (x"49",x"87",x"eb",x"c2"),
  1451 => (x"69",x"97",x"81",x"cb"),
  1452 => (x"02",x"99",x"d0",x"49"),
  1453 => (x"c1",x"87",x"d9",x"c1"),
  1454 => (x"74",x"4b",x"d0",x"d6"),
  1455 => (x"c1",x"91",x"cc",x"49"),
  1456 => (x"c8",x"81",x"c4",x"f7"),
  1457 => (x"7a",x"73",x"4a",x"a1"),
  1458 => (x"ff",x"c3",x"81",x"c1"),
  1459 => (x"de",x"49",x"74",x"51"),
  1460 => (x"d8",x"fb",x"c2",x"91"),
  1461 => (x"c2",x"85",x"71",x"4d"),
  1462 => (x"c1",x"7d",x"97",x"c1"),
  1463 => (x"e0",x"c0",x"49",x"a5"),
  1464 => (x"e8",x"f5",x"c2",x"51"),
  1465 => (x"d2",x"02",x"bf",x"97"),
  1466 => (x"c2",x"84",x"c1",x"87"),
  1467 => (x"f5",x"c2",x"4b",x"a5"),
  1468 => (x"49",x"db",x"4a",x"e8"),
  1469 => (x"87",x"d3",x"eb",x"fe"),
  1470 => (x"cd",x"87",x"db",x"c1"),
  1471 => (x"51",x"c0",x"49",x"a5"),
  1472 => (x"a5",x"c2",x"84",x"c1"),
  1473 => (x"cb",x"4a",x"6e",x"4b"),
  1474 => (x"fe",x"ea",x"fe",x"49"),
  1475 => (x"87",x"c6",x"c1",x"87"),
  1476 => (x"91",x"cc",x"49",x"74"),
  1477 => (x"81",x"c4",x"f7",x"c1"),
  1478 => (x"d4",x"c1",x"81",x"c8"),
  1479 => (x"f5",x"c2",x"79",x"df"),
  1480 => (x"02",x"bf",x"97",x"e8"),
  1481 => (x"49",x"74",x"87",x"d8"),
  1482 => (x"84",x"c1",x"91",x"de"),
  1483 => (x"4b",x"d8",x"fb",x"c2"),
  1484 => (x"f5",x"c2",x"83",x"71"),
  1485 => (x"49",x"dd",x"4a",x"e8"),
  1486 => (x"87",x"cf",x"ea",x"fe"),
  1487 => (x"4b",x"74",x"87",x"d8"),
  1488 => (x"fb",x"c2",x"93",x"de"),
  1489 => (x"a3",x"cb",x"83",x"d8"),
  1490 => (x"c1",x"51",x"c0",x"49"),
  1491 => (x"4a",x"6e",x"73",x"84"),
  1492 => (x"e9",x"fe",x"49",x"cb"),
  1493 => (x"66",x"c4",x"87",x"f5"),
  1494 => (x"c8",x"80",x"c1",x"48"),
  1495 => (x"b7",x"c7",x"58",x"a6"),
  1496 => (x"c5",x"c0",x"03",x"ac"),
  1497 => (x"fc",x"05",x"6e",x"87"),
  1498 => (x"b7",x"c7",x"87",x"dd"),
  1499 => (x"d3",x"c0",x"03",x"ac"),
  1500 => (x"de",x"49",x"74",x"87"),
  1501 => (x"d8",x"fb",x"c2",x"91"),
  1502 => (x"c1",x"51",x"c0",x"81"),
  1503 => (x"ac",x"b7",x"c7",x"84"),
  1504 => (x"87",x"ed",x"ff",x"04"),
  1505 => (x"48",x"d9",x"f8",x"c1"),
  1506 => (x"f8",x"c1",x"50",x"c0"),
  1507 => (x"50",x"c2",x"48",x"d8"),
  1508 => (x"48",x"e0",x"f8",x"c1"),
  1509 => (x"78",x"c2",x"df",x"c1"),
  1510 => (x"48",x"dc",x"f8",x"c1"),
  1511 => (x"78",x"d2",x"d2",x"c1"),
  1512 => (x"48",x"ec",x"f8",x"c1"),
  1513 => (x"78",x"f6",x"d6",x"c1"),
  1514 => (x"c0",x"49",x"66",x"cc"),
  1515 => (x"f0",x"87",x"f3",x"fb"),
  1516 => (x"87",x"db",x"e6",x"8e"),
  1517 => (x"c2",x"4a",x"71",x"1e"),
  1518 => (x"72",x"5a",x"f4",x"fa"),
  1519 => (x"87",x"dc",x"f9",x"49"),
  1520 => (x"71",x"1e",x"4f",x"26"),
  1521 => (x"91",x"cc",x"49",x"4a"),
  1522 => (x"81",x"c4",x"f7",x"c1"),
  1523 => (x"48",x"11",x"81",x"c1"),
  1524 => (x"58",x"f0",x"fa",x"c2"),
  1525 => (x"49",x"a2",x"f0",x"c0"),
  1526 => (x"87",x"ff",x"e7",x"fe"),
  1527 => (x"dd",x"d5",x"49",x"c0"),
  1528 => (x"0e",x"4f",x"26",x"87"),
  1529 => (x"5d",x"5c",x"5b",x"5e"),
  1530 => (x"71",x"86",x"f0",x"0e"),
  1531 => (x"91",x"cc",x"49",x"4c"),
  1532 => (x"81",x"c4",x"f7",x"c1"),
  1533 => (x"c4",x"7e",x"a1",x"c3"),
  1534 => (x"fa",x"c2",x"48",x"a6"),
  1535 => (x"6e",x"78",x"bf",x"e8"),
  1536 => (x"c4",x"4a",x"bf",x"97"),
  1537 => (x"2b",x"72",x"4b",x"66"),
  1538 => (x"12",x"4a",x"a1",x"c1"),
  1539 => (x"58",x"a6",x"cc",x"48"),
  1540 => (x"83",x"c1",x"9b",x"70"),
  1541 => (x"69",x"97",x"81",x"c2"),
  1542 => (x"04",x"ab",x"b7",x"49"),
  1543 => (x"4b",x"c0",x"87",x"c2"),
  1544 => (x"4a",x"bf",x"97",x"6e"),
  1545 => (x"72",x"49",x"66",x"c8"),
  1546 => (x"c4",x"b9",x"ff",x"31"),
  1547 => (x"4d",x"73",x"99",x"66"),
  1548 => (x"b5",x"71",x"35",x"72"),
  1549 => (x"5d",x"ec",x"fa",x"c2"),
  1550 => (x"c3",x"48",x"d4",x"ff"),
  1551 => (x"d0",x"ff",x"78",x"ff"),
  1552 => (x"c0",x"c8",x"48",x"bf"),
  1553 => (x"a6",x"d0",x"98",x"c0"),
  1554 => (x"02",x"98",x"70",x"58"),
  1555 => (x"d0",x"ff",x"87",x"d0"),
  1556 => (x"c0",x"c8",x"48",x"bf"),
  1557 => (x"a6",x"c4",x"98",x"c0"),
  1558 => (x"05",x"98",x"70",x"58"),
  1559 => (x"d0",x"ff",x"87",x"f0"),
  1560 => (x"78",x"e1",x"c0",x"48"),
  1561 => (x"de",x"48",x"d4",x"ff"),
  1562 => (x"7d",x"0d",x"70",x"78"),
  1563 => (x"c8",x"48",x"75",x"0d"),
  1564 => (x"d4",x"ff",x"28",x"b7"),
  1565 => (x"48",x"75",x"78",x"08"),
  1566 => (x"ff",x"28",x"b7",x"d0"),
  1567 => (x"75",x"78",x"08",x"d4"),
  1568 => (x"28",x"b7",x"d8",x"48"),
  1569 => (x"78",x"08",x"d4",x"ff"),
  1570 => (x"48",x"bf",x"d0",x"ff"),
  1571 => (x"98",x"c0",x"c0",x"c8"),
  1572 => (x"70",x"58",x"a6",x"c4"),
  1573 => (x"87",x"d0",x"02",x"98"),
  1574 => (x"48",x"bf",x"d0",x"ff"),
  1575 => (x"98",x"c0",x"c0",x"c8"),
  1576 => (x"70",x"58",x"a6",x"c4"),
  1577 => (x"87",x"f0",x"05",x"98"),
  1578 => (x"c0",x"48",x"d0",x"ff"),
  1579 => (x"1e",x"c7",x"78",x"e0"),
  1580 => (x"f7",x"c1",x"1e",x"c0"),
  1581 => (x"fa",x"c2",x"1e",x"c4"),
  1582 => (x"c1",x"49",x"bf",x"ec"),
  1583 => (x"49",x"74",x"87",x"e1"),
  1584 => (x"87",x"de",x"f7",x"c0"),
  1585 => (x"c6",x"e2",x"8e",x"e4"),
  1586 => (x"1e",x"73",x"1e",x"87"),
  1587 => (x"fc",x"49",x"4b",x"71"),
  1588 => (x"49",x"73",x"87",x"d1"),
  1589 => (x"e1",x"87",x"cc",x"fc"),
  1590 => (x"73",x"1e",x"87",x"f9"),
  1591 => (x"c2",x"4b",x"71",x"1e"),
  1592 => (x"d5",x"02",x"4a",x"a3"),
  1593 => (x"05",x"8a",x"c1",x"87"),
  1594 => (x"fb",x"c2",x"87",x"db"),
  1595 => (x"d4",x"02",x"bf",x"c0"),
  1596 => (x"88",x"c1",x"48",x"87"),
  1597 => (x"58",x"c4",x"fb",x"c2"),
  1598 => (x"fb",x"c2",x"87",x"cb"),
  1599 => (x"c1",x"48",x"bf",x"c0"),
  1600 => (x"c4",x"fb",x"c2",x"80"),
  1601 => (x"c0",x"1e",x"c7",x"58"),
  1602 => (x"c4",x"f7",x"c1",x"1e"),
  1603 => (x"ec",x"fa",x"c2",x"1e"),
  1604 => (x"87",x"cb",x"49",x"bf"),
  1605 => (x"f6",x"c0",x"49",x"73"),
  1606 => (x"8e",x"f4",x"87",x"c8"),
  1607 => (x"0e",x"87",x"f4",x"e0"),
  1608 => (x"5d",x"5c",x"5b",x"5e"),
  1609 => (x"86",x"d8",x"ff",x"0e"),
  1610 => (x"c8",x"59",x"a6",x"dc"),
  1611 => (x"78",x"c0",x"48",x"a6"),
  1612 => (x"78",x"c0",x"80",x"c4"),
  1613 => (x"c2",x"80",x"c4",x"4d"),
  1614 => (x"78",x"bf",x"c0",x"fb"),
  1615 => (x"c3",x"48",x"d4",x"ff"),
  1616 => (x"d0",x"ff",x"78",x"ff"),
  1617 => (x"c0",x"c8",x"48",x"bf"),
  1618 => (x"a6",x"c4",x"98",x"c0"),
  1619 => (x"02",x"98",x"70",x"58"),
  1620 => (x"d0",x"ff",x"87",x"d0"),
  1621 => (x"c0",x"c8",x"48",x"bf"),
  1622 => (x"a6",x"c4",x"98",x"c0"),
  1623 => (x"05",x"98",x"70",x"58"),
  1624 => (x"d0",x"ff",x"87",x"f0"),
  1625 => (x"78",x"e1",x"c0",x"48"),
  1626 => (x"d4",x"48",x"d4",x"ff"),
  1627 => (x"d5",x"dd",x"ff",x"78"),
  1628 => (x"48",x"d4",x"ff",x"87"),
  1629 => (x"d4",x"78",x"ff",x"c3"),
  1630 => (x"d4",x"ff",x"48",x"a6"),
  1631 => (x"66",x"d4",x"78",x"bf"),
  1632 => (x"a8",x"fb",x"c0",x"48"),
  1633 => (x"87",x"d3",x"c1",x"02"),
  1634 => (x"4a",x"66",x"f8",x"c0"),
  1635 => (x"7e",x"6a",x"82",x"c4"),
  1636 => (x"d2",x"c1",x"1e",x"72"),
  1637 => (x"66",x"c4",x"48",x"d9"),
  1638 => (x"4a",x"a1",x"c8",x"49"),
  1639 => (x"aa",x"71",x"41",x"20"),
  1640 => (x"10",x"87",x"f9",x"05"),
  1641 => (x"c0",x"4a",x"26",x"51"),
  1642 => (x"c8",x"49",x"66",x"f8"),
  1643 => (x"f4",x"de",x"c1",x"81"),
  1644 => (x"c7",x"49",x"6a",x"79"),
  1645 => (x"51",x"66",x"d4",x"81"),
  1646 => (x"1e",x"d8",x"1e",x"c1"),
  1647 => (x"81",x"c8",x"49",x"6a"),
  1648 => (x"87",x"d9",x"dc",x"ff"),
  1649 => (x"66",x"d0",x"86",x"c8"),
  1650 => (x"a8",x"b7",x"c0",x"48"),
  1651 => (x"c1",x"87",x"c4",x"01"),
  1652 => (x"d0",x"87",x"c8",x"4d"),
  1653 => (x"88",x"c1",x"48",x"66"),
  1654 => (x"d4",x"58",x"a6",x"d4"),
  1655 => (x"f4",x"ca",x"02",x"66"),
  1656 => (x"66",x"c0",x"c1",x"87"),
  1657 => (x"ca",x"03",x"ad",x"b7"),
  1658 => (x"d4",x"ff",x"87",x"eb"),
  1659 => (x"78",x"ff",x"c3",x"48"),
  1660 => (x"ff",x"48",x"a6",x"d4"),
  1661 => (x"d4",x"78",x"bf",x"d4"),
  1662 => (x"c6",x"c1",x"48",x"66"),
  1663 => (x"58",x"a6",x"c4",x"88"),
  1664 => (x"c0",x"02",x"98",x"70"),
  1665 => (x"c9",x"48",x"87",x"e6"),
  1666 => (x"58",x"a6",x"c4",x"88"),
  1667 => (x"c4",x"02",x"98",x"70"),
  1668 => (x"c1",x"48",x"87",x"d5"),
  1669 => (x"58",x"a6",x"c4",x"88"),
  1670 => (x"c1",x"02",x"98",x"70"),
  1671 => (x"c4",x"48",x"87",x"e3"),
  1672 => (x"70",x"58",x"a6",x"88"),
  1673 => (x"fe",x"c3",x"02",x"98"),
  1674 => (x"87",x"d3",x"c9",x"87"),
  1675 => (x"c1",x"05",x"66",x"d8"),
  1676 => (x"d4",x"ff",x"87",x"c5"),
  1677 => (x"78",x"ff",x"c3",x"48"),
  1678 => (x"1e",x"ca",x"1e",x"c0"),
  1679 => (x"93",x"cc",x"4b",x"75"),
  1680 => (x"83",x"66",x"c0",x"c1"),
  1681 => (x"6c",x"4c",x"a3",x"c4"),
  1682 => (x"d0",x"da",x"ff",x"49"),
  1683 => (x"de",x"1e",x"c1",x"87"),
  1684 => (x"ff",x"49",x"6c",x"1e"),
  1685 => (x"d0",x"87",x"c6",x"da"),
  1686 => (x"49",x"a3",x"c8",x"86"),
  1687 => (x"79",x"f4",x"de",x"c1"),
  1688 => (x"ad",x"b7",x"66",x"d0"),
  1689 => (x"c1",x"87",x"c5",x"04"),
  1690 => (x"87",x"da",x"c8",x"85"),
  1691 => (x"c1",x"48",x"66",x"d0"),
  1692 => (x"58",x"a6",x"d4",x"88"),
  1693 => (x"ff",x"87",x"cf",x"c8"),
  1694 => (x"d8",x"87",x"cb",x"d9"),
  1695 => (x"c5",x"c8",x"58",x"a6"),
  1696 => (x"d2",x"db",x"ff",x"87"),
  1697 => (x"58",x"a6",x"cc",x"87"),
  1698 => (x"a8",x"b7",x"66",x"cc"),
  1699 => (x"cc",x"87",x"c6",x"06"),
  1700 => (x"66",x"c8",x"48",x"a6"),
  1701 => (x"fe",x"da",x"ff",x"78"),
  1702 => (x"a8",x"ec",x"c0",x"87"),
  1703 => (x"87",x"c7",x"c2",x"05"),
  1704 => (x"c1",x"05",x"66",x"d8"),
  1705 => (x"49",x"75",x"87",x"f7"),
  1706 => (x"f8",x"c0",x"91",x"cc"),
  1707 => (x"a1",x"c4",x"81",x"66"),
  1708 => (x"c1",x"4c",x"6a",x"4a"),
  1709 => (x"66",x"c8",x"4a",x"a1"),
  1710 => (x"79",x"97",x"c2",x"52"),
  1711 => (x"df",x"c1",x"81",x"c8"),
  1712 => (x"d4",x"ff",x"79",x"c2"),
  1713 => (x"78",x"ff",x"c3",x"48"),
  1714 => (x"ff",x"48",x"a6",x"d4"),
  1715 => (x"d4",x"78",x"bf",x"d4"),
  1716 => (x"e8",x"c0",x"02",x"66"),
  1717 => (x"fb",x"c0",x"48",x"87"),
  1718 => (x"e0",x"c0",x"02",x"a8"),
  1719 => (x"97",x"66",x"d4",x"87"),
  1720 => (x"ff",x"84",x"c1",x"7c"),
  1721 => (x"ff",x"c3",x"48",x"d4"),
  1722 => (x"48",x"a6",x"d4",x"78"),
  1723 => (x"78",x"bf",x"d4",x"ff"),
  1724 => (x"c8",x"02",x"66",x"d4"),
  1725 => (x"fb",x"c0",x"48",x"87"),
  1726 => (x"e0",x"ff",x"05",x"a8"),
  1727 => (x"54",x"e0",x"c0",x"87"),
  1728 => (x"c0",x"54",x"c1",x"c2"),
  1729 => (x"66",x"d0",x"7c",x"97"),
  1730 => (x"c5",x"04",x"ad",x"b7"),
  1731 => (x"c5",x"85",x"c1",x"87"),
  1732 => (x"66",x"d0",x"87",x"f4"),
  1733 => (x"d4",x"88",x"c1",x"48"),
  1734 => (x"e9",x"c5",x"58",x"a6"),
  1735 => (x"e5",x"d6",x"ff",x"87"),
  1736 => (x"58",x"a6",x"d8",x"87"),
  1737 => (x"c8",x"87",x"df",x"c5"),
  1738 => (x"66",x"d8",x"48",x"66"),
  1739 => (x"c4",x"c5",x"05",x"a8"),
  1740 => (x"48",x"a6",x"dc",x"87"),
  1741 => (x"d8",x"ff",x"78",x"c0"),
  1742 => (x"a6",x"d8",x"87",x"dd"),
  1743 => (x"d6",x"d8",x"ff",x"58"),
  1744 => (x"a6",x"e4",x"c0",x"87"),
  1745 => (x"a8",x"ec",x"c0",x"58"),
  1746 => (x"87",x"ca",x"c0",x"05"),
  1747 => (x"48",x"a6",x"e0",x"c0"),
  1748 => (x"c0",x"78",x"66",x"d4"),
  1749 => (x"d4",x"ff",x"87",x"c6"),
  1750 => (x"78",x"ff",x"c3",x"48"),
  1751 => (x"91",x"cc",x"49",x"75"),
  1752 => (x"48",x"66",x"f8",x"c0"),
  1753 => (x"a6",x"c4",x"80",x"71"),
  1754 => (x"c3",x"49",x"6e",x"58"),
  1755 => (x"51",x"66",x"d4",x"81"),
  1756 => (x"49",x"66",x"e0",x"c0"),
  1757 => (x"66",x"d4",x"81",x"c1"),
  1758 => (x"71",x"48",x"c1",x"89"),
  1759 => (x"c1",x"49",x"70",x"30"),
  1760 => (x"c1",x"4a",x"6e",x"89"),
  1761 => (x"97",x"09",x"72",x"82"),
  1762 => (x"48",x"6e",x"09",x"79"),
  1763 => (x"fa",x"c2",x"50",x"c2"),
  1764 => (x"d4",x"49",x"bf",x"e8"),
  1765 => (x"97",x"29",x"b7",x"66"),
  1766 => (x"71",x"48",x"4a",x"6a"),
  1767 => (x"a6",x"e8",x"c0",x"98"),
  1768 => (x"c4",x"48",x"6e",x"58"),
  1769 => (x"58",x"a6",x"c8",x"80"),
  1770 => (x"4c",x"bf",x"66",x"c4"),
  1771 => (x"c8",x"48",x"66",x"d8"),
  1772 => (x"c0",x"02",x"a8",x"66"),
  1773 => (x"e0",x"c0",x"87",x"c9"),
  1774 => (x"78",x"c0",x"48",x"a6"),
  1775 => (x"c0",x"87",x"c6",x"c0"),
  1776 => (x"c1",x"48",x"a6",x"e0"),
  1777 => (x"66",x"e0",x"c0",x"78"),
  1778 => (x"1e",x"e0",x"c0",x"1e"),
  1779 => (x"d4",x"ff",x"49",x"74"),
  1780 => (x"86",x"c8",x"87",x"cb"),
  1781 => (x"c0",x"58",x"a6",x"d8"),
  1782 => (x"c1",x"06",x"a8",x"b7"),
  1783 => (x"66",x"d4",x"87",x"da"),
  1784 => (x"bf",x"66",x"c4",x"84"),
  1785 => (x"81",x"e0",x"c0",x"49"),
  1786 => (x"c1",x"4b",x"89",x"74"),
  1787 => (x"71",x"4a",x"e2",x"d2"),
  1788 => (x"87",x"d7",x"d7",x"fe"),
  1789 => (x"66",x"dc",x"84",x"c2"),
  1790 => (x"c0",x"80",x"c1",x"48"),
  1791 => (x"c0",x"58",x"a6",x"e0"),
  1792 => (x"c1",x"49",x"66",x"e4"),
  1793 => (x"02",x"a9",x"70",x"81"),
  1794 => (x"c0",x"87",x"c9",x"c0"),
  1795 => (x"c0",x"48",x"a6",x"e0"),
  1796 => (x"87",x"c6",x"c0",x"78"),
  1797 => (x"48",x"a6",x"e0",x"c0"),
  1798 => (x"e0",x"c0",x"78",x"c1"),
  1799 => (x"66",x"c8",x"1e",x"66"),
  1800 => (x"e0",x"c0",x"49",x"bf"),
  1801 => (x"71",x"89",x"74",x"81"),
  1802 => (x"ff",x"49",x"74",x"1e"),
  1803 => (x"c8",x"87",x"ee",x"d2"),
  1804 => (x"a8",x"b7",x"c0",x"86"),
  1805 => (x"87",x"fe",x"fe",x"01"),
  1806 => (x"c0",x"02",x"66",x"dc"),
  1807 => (x"49",x"6e",x"87",x"d2"),
  1808 => (x"66",x"dc",x"81",x"c2"),
  1809 => (x"c8",x"49",x"6e",x"51"),
  1810 => (x"e3",x"df",x"c1",x"81"),
  1811 => (x"87",x"cd",x"c0",x"79"),
  1812 => (x"81",x"c2",x"49",x"6e"),
  1813 => (x"c8",x"49",x"6e",x"51"),
  1814 => (x"c9",x"e3",x"c1",x"81"),
  1815 => (x"b7",x"66",x"d0",x"79"),
  1816 => (x"c5",x"c0",x"04",x"ad"),
  1817 => (x"c0",x"85",x"c1",x"87"),
  1818 => (x"66",x"d0",x"87",x"dc"),
  1819 => (x"d4",x"88",x"c1",x"48"),
  1820 => (x"d1",x"c0",x"58",x"a6"),
  1821 => (x"cd",x"d1",x"ff",x"87"),
  1822 => (x"58",x"a6",x"d8",x"87"),
  1823 => (x"ff",x"87",x"c7",x"c0"),
  1824 => (x"d8",x"87",x"c3",x"d1"),
  1825 => (x"66",x"d4",x"58",x"a6"),
  1826 => (x"87",x"c9",x"c0",x"02"),
  1827 => (x"b7",x"66",x"c0",x"c1"),
  1828 => (x"d5",x"f5",x"04",x"ad"),
  1829 => (x"ad",x"b7",x"c7",x"87"),
  1830 => (x"87",x"dc",x"c0",x"03"),
  1831 => (x"91",x"cc",x"49",x"75"),
  1832 => (x"81",x"66",x"f8",x"c0"),
  1833 => (x"6a",x"4a",x"a1",x"c4"),
  1834 => (x"c8",x"52",x"c0",x"4a"),
  1835 => (x"c1",x"79",x"c0",x"81"),
  1836 => (x"ad",x"b7",x"c7",x"85"),
  1837 => (x"87",x"e4",x"ff",x"04"),
  1838 => (x"c0",x"02",x"66",x"d8"),
  1839 => (x"f8",x"c0",x"87",x"eb"),
  1840 => (x"d4",x"c1",x"49",x"66"),
  1841 => (x"66",x"f8",x"c0",x"81"),
  1842 => (x"82",x"d5",x"c1",x"4a"),
  1843 => (x"51",x"c2",x"52",x"c0"),
  1844 => (x"49",x"66",x"f8",x"c0"),
  1845 => (x"c1",x"81",x"dc",x"c1"),
  1846 => (x"c0",x"79",x"c2",x"df"),
  1847 => (x"c1",x"49",x"66",x"f8"),
  1848 => (x"d2",x"c1",x"81",x"d8"),
  1849 => (x"d6",x"c0",x"79",x"e5"),
  1850 => (x"66",x"f8",x"c0",x"87"),
  1851 => (x"81",x"d8",x"c1",x"49"),
  1852 => (x"79",x"ec",x"d2",x"c1"),
  1853 => (x"49",x"66",x"f8",x"c0"),
  1854 => (x"c2",x"81",x"dc",x"c1"),
  1855 => (x"c1",x"79",x"cd",x"de"),
  1856 => (x"c0",x"4a",x"da",x"e3"),
  1857 => (x"c1",x"49",x"66",x"f8"),
  1858 => (x"79",x"72",x"81",x"e8"),
  1859 => (x"48",x"bf",x"d0",x"ff"),
  1860 => (x"98",x"c0",x"c0",x"c8"),
  1861 => (x"70",x"58",x"a6",x"c4"),
  1862 => (x"d1",x"c0",x"02",x"98"),
  1863 => (x"bf",x"d0",x"ff",x"87"),
  1864 => (x"c0",x"c0",x"c8",x"48"),
  1865 => (x"58",x"a6",x"c4",x"98"),
  1866 => (x"ff",x"05",x"98",x"70"),
  1867 => (x"d0",x"ff",x"87",x"ef"),
  1868 => (x"78",x"e0",x"c0",x"48"),
  1869 => (x"ff",x"48",x"66",x"cc"),
  1870 => (x"d0",x"ff",x"8e",x"d8"),
  1871 => (x"c7",x"1e",x"87",x"d1"),
  1872 => (x"c1",x"1e",x"c0",x"1e"),
  1873 => (x"c2",x"1e",x"c4",x"f7"),
  1874 => (x"49",x"bf",x"ec",x"fa"),
  1875 => (x"c1",x"87",x"d0",x"ef"),
  1876 => (x"c0",x"49",x"c4",x"f7"),
  1877 => (x"f4",x"87",x"d6",x"e8"),
  1878 => (x"1e",x"4f",x"26",x"8e"),
  1879 => (x"c2",x"87",x"c6",x"ca"),
  1880 => (x"c0",x"48",x"c8",x"fb"),
  1881 => (x"48",x"d4",x"ff",x"50"),
  1882 => (x"c1",x"78",x"ff",x"c3"),
  1883 => (x"fe",x"49",x"f3",x"d2"),
  1884 => (x"fe",x"87",x"f4",x"d0"),
  1885 => (x"70",x"87",x"f0",x"dd"),
  1886 => (x"87",x"cd",x"02",x"98"),
  1887 => (x"87",x"f0",x"ea",x"fe"),
  1888 => (x"c4",x"02",x"98",x"70"),
  1889 => (x"c2",x"4a",x"c1",x"87"),
  1890 => (x"72",x"4a",x"c0",x"87"),
  1891 => (x"87",x"c8",x"02",x"9a"),
  1892 => (x"49",x"c9",x"d3",x"c1"),
  1893 => (x"87",x"cf",x"d0",x"fe"),
  1894 => (x"bf",x"d8",x"ec",x"c2"),
  1895 => (x"c2",x"d4",x"ff",x"49"),
  1896 => (x"c0",x"fb",x"c2",x"87"),
  1897 => (x"c2",x"78",x"c0",x"48"),
  1898 => (x"c0",x"48",x"ec",x"fa"),
  1899 => (x"cd",x"fe",x"49",x"78"),
  1900 => (x"87",x"dd",x"c3",x"87"),
  1901 => (x"c0",x"87",x"c2",x"c9"),
  1902 => (x"ff",x"87",x"e1",x"e7"),
  1903 => (x"4f",x"26",x"87",x"f6"),
  1904 => (x"00",x"00",x"14",x"d2"),
  1905 => (x"00",x"00",x"00",x"02"),
  1906 => (x"00",x"00",x"2e",x"d8"),
  1907 => (x"00",x"00",x"15",x"1f"),
  1908 => (x"00",x"00",x"00",x"02"),
  1909 => (x"00",x"00",x"2e",x"f6"),
  1910 => (x"00",x"00",x"15",x"1f"),
  1911 => (x"00",x"00",x"00",x"02"),
  1912 => (x"00",x"00",x"2f",x"14"),
  1913 => (x"00",x"00",x"15",x"1f"),
  1914 => (x"00",x"00",x"00",x"02"),
  1915 => (x"00",x"00",x"2f",x"32"),
  1916 => (x"00",x"00",x"15",x"1f"),
  1917 => (x"00",x"00",x"00",x"02"),
  1918 => (x"00",x"00",x"2f",x"50"),
  1919 => (x"00",x"00",x"15",x"1f"),
  1920 => (x"00",x"00",x"00",x"02"),
  1921 => (x"00",x"00",x"2f",x"6e"),
  1922 => (x"00",x"00",x"15",x"1f"),
  1923 => (x"00",x"00",x"00",x"02"),
  1924 => (x"00",x"00",x"2f",x"8c"),
  1925 => (x"00",x"00",x"15",x"1f"),
  1926 => (x"00",x"00",x"00",x"02"),
  1927 => (x"00",x"00",x"00",x"00"),
  1928 => (x"00",x"00",x"17",x"c2"),
  1929 => (x"00",x"00",x"00",x"00"),
  1930 => (x"00",x"00",x"00",x"00"),
  1931 => (x"00",x"00",x"15",x"b6"),
  1932 => (x"d5",x"c1",x"1e",x"1e"),
  1933 => (x"58",x"a6",x"c4",x"87"),
  1934 => (x"1e",x"4f",x"26",x"26"),
  1935 => (x"f0",x"fe",x"4a",x"71"),
  1936 => (x"cd",x"78",x"c0",x"48"),
  1937 => (x"c1",x"0a",x"7a",x"0a"),
  1938 => (x"fe",x"49",x"d1",x"f9"),
  1939 => (x"26",x"87",x"d8",x"cd"),
  1940 => (x"74",x"65",x"53",x"4f"),
  1941 => (x"6e",x"61",x"68",x"20"),
  1942 => (x"72",x"65",x"6c",x"64"),
  1943 => (x"6e",x"49",x"00",x"0a"),
  1944 => (x"74",x"6e",x"69",x"20"),
  1945 => (x"75",x"72",x"72",x"65"),
  1946 => (x"63",x"20",x"74",x"70"),
  1947 => (x"74",x"73",x"6e",x"6f"),
  1948 => (x"74",x"63",x"75",x"72"),
  1949 => (x"00",x"0a",x"72",x"6f"),
  1950 => (x"de",x"f9",x"c1",x"1e"),
  1951 => (x"e6",x"cc",x"fe",x"49"),
  1952 => (x"f0",x"f8",x"c1",x"87"),
  1953 => (x"87",x"f3",x"fe",x"49"),
  1954 => (x"fe",x"1e",x"4f",x"26"),
  1955 => (x"26",x"48",x"bf",x"f0"),
  1956 => (x"f0",x"fe",x"1e",x"4f"),
  1957 => (x"26",x"78",x"c1",x"48"),
  1958 => (x"f0",x"fe",x"1e",x"4f"),
  1959 => (x"26",x"78",x"c0",x"48"),
  1960 => (x"4a",x"71",x"1e",x"4f"),
  1961 => (x"a2",x"c4",x"7a",x"c0"),
  1962 => (x"c8",x"79",x"c0",x"49"),
  1963 => (x"79",x"c0",x"49",x"a2"),
  1964 => (x"c0",x"49",x"a2",x"cc"),
  1965 => (x"0e",x"4f",x"26",x"79"),
  1966 => (x"0e",x"5c",x"5b",x"5e"),
  1967 => (x"4c",x"71",x"86",x"f8"),
  1968 => (x"cc",x"49",x"a4",x"c8"),
  1969 => (x"48",x"6b",x"4b",x"a4"),
  1970 => (x"a6",x"c4",x"80",x"c1"),
  1971 => (x"c8",x"98",x"cf",x"58"),
  1972 => (x"48",x"69",x"58",x"a6"),
  1973 => (x"05",x"a8",x"66",x"c4"),
  1974 => (x"48",x"6b",x"87",x"d4"),
  1975 => (x"a6",x"c4",x"80",x"c1"),
  1976 => (x"c8",x"98",x"cf",x"58"),
  1977 => (x"48",x"69",x"58",x"a6"),
  1978 => (x"02",x"a8",x"66",x"c4"),
  1979 => (x"e8",x"fe",x"87",x"ec"),
  1980 => (x"a4",x"d0",x"c1",x"87"),
  1981 => (x"c4",x"48",x"6b",x"49"),
  1982 => (x"58",x"a6",x"c4",x"90"),
  1983 => (x"66",x"d4",x"81",x"70"),
  1984 => (x"c1",x"48",x"6b",x"79"),
  1985 => (x"58",x"a6",x"c8",x"80"),
  1986 => (x"7b",x"70",x"98",x"cf"),
  1987 => (x"fd",x"87",x"d2",x"c1"),
  1988 => (x"8e",x"f8",x"87",x"ff"),
  1989 => (x"4d",x"26",x"87",x"c2"),
  1990 => (x"4b",x"26",x"4c",x"26"),
  1991 => (x"5e",x"0e",x"4f",x"26"),
  1992 => (x"0e",x"5d",x"5c",x"5b"),
  1993 => (x"4d",x"71",x"86",x"f8"),
  1994 => (x"6d",x"4c",x"a5",x"c4"),
  1995 => (x"05",x"a8",x"6c",x"48"),
  1996 => (x"48",x"ff",x"87",x"c5"),
  1997 => (x"fd",x"87",x"e5",x"c0"),
  1998 => (x"a5",x"d0",x"87",x"df"),
  1999 => (x"c4",x"48",x"6c",x"4b"),
  2000 => (x"58",x"a6",x"c4",x"90"),
  2001 => (x"4b",x"6b",x"83",x"70"),
  2002 => (x"6c",x"9b",x"ff",x"c3"),
  2003 => (x"c8",x"80",x"c1",x"48"),
  2004 => (x"98",x"cf",x"58",x"a6"),
  2005 => (x"f8",x"fc",x"7c",x"70"),
  2006 => (x"48",x"49",x"73",x"87"),
  2007 => (x"f5",x"fe",x"8e",x"f8"),
  2008 => (x"1e",x"73",x"1e",x"87"),
  2009 => (x"f0",x"fc",x"86",x"f8"),
  2010 => (x"4b",x"bf",x"e0",x"87"),
  2011 => (x"c0",x"e0",x"c0",x"49"),
  2012 => (x"e7",x"c0",x"02",x"99"),
  2013 => (x"c3",x"4a",x"73",x"87"),
  2014 => (x"fe",x"c2",x"9a",x"ff"),
  2015 => (x"c4",x"48",x"bf",x"ea"),
  2016 => (x"58",x"a6",x"c4",x"90"),
  2017 => (x"49",x"fa",x"fe",x"c2"),
  2018 => (x"79",x"72",x"81",x"70"),
  2019 => (x"bf",x"ea",x"fe",x"c2"),
  2020 => (x"c8",x"80",x"c1",x"48"),
  2021 => (x"98",x"cf",x"58",x"a6"),
  2022 => (x"58",x"ee",x"fe",x"c2"),
  2023 => (x"c0",x"d0",x"49",x"73"),
  2024 => (x"f2",x"c0",x"02",x"99"),
  2025 => (x"f2",x"fe",x"c2",x"87"),
  2026 => (x"fe",x"c2",x"48",x"bf"),
  2027 => (x"02",x"a8",x"bf",x"f6"),
  2028 => (x"c2",x"87",x"e4",x"c0"),
  2029 => (x"48",x"bf",x"f2",x"fe"),
  2030 => (x"a6",x"c4",x"90",x"c4"),
  2031 => (x"fa",x"ff",x"c2",x"58"),
  2032 => (x"e0",x"81",x"70",x"49"),
  2033 => (x"c2",x"78",x"69",x"48"),
  2034 => (x"48",x"bf",x"f2",x"fe"),
  2035 => (x"a6",x"c8",x"80",x"c1"),
  2036 => (x"c2",x"98",x"cf",x"58"),
  2037 => (x"fa",x"58",x"f6",x"fe"),
  2038 => (x"a6",x"c4",x"87",x"f0"),
  2039 => (x"87",x"f1",x"fa",x"58"),
  2040 => (x"f5",x"fc",x"8e",x"f8"),
  2041 => (x"fe",x"c2",x"1e",x"87"),
  2042 => (x"f4",x"fa",x"49",x"ea"),
  2043 => (x"e1",x"fd",x"c1",x"87"),
  2044 => (x"87",x"c7",x"f9",x"49"),
  2045 => (x"26",x"87",x"f5",x"c3"),
  2046 => (x"1e",x"73",x"1e",x"4f"),
  2047 => (x"49",x"ea",x"fe",x"c2"),
  2048 => (x"70",x"87",x"db",x"fc"),
  2049 => (x"aa",x"b7",x"c0",x"4a"),
  2050 => (x"87",x"cc",x"c2",x"04"),
  2051 => (x"05",x"aa",x"f0",x"c3"),
  2052 => (x"c2",x"c2",x"87",x"c9"),
  2053 => (x"78",x"c1",x"48",x"e4"),
  2054 => (x"c3",x"87",x"ed",x"c1"),
  2055 => (x"c9",x"05",x"aa",x"e0"),
  2056 => (x"e8",x"c2",x"c2",x"87"),
  2057 => (x"c1",x"78",x"c1",x"48"),
  2058 => (x"c2",x"c2",x"87",x"de"),
  2059 => (x"c6",x"02",x"bf",x"e8"),
  2060 => (x"a2",x"c0",x"c2",x"87"),
  2061 => (x"72",x"87",x"c2",x"4b"),
  2062 => (x"e4",x"c2",x"c2",x"4b"),
  2063 => (x"e0",x"c0",x"02",x"bf"),
  2064 => (x"c4",x"49",x"73",x"87"),
  2065 => (x"c2",x"91",x"29",x"b7"),
  2066 => (x"73",x"81",x"ec",x"c2"),
  2067 => (x"c2",x"9a",x"cf",x"4a"),
  2068 => (x"72",x"48",x"c1",x"92"),
  2069 => (x"ff",x"4a",x"70",x"30"),
  2070 => (x"69",x"48",x"72",x"ba"),
  2071 => (x"db",x"79",x"70",x"98"),
  2072 => (x"c4",x"49",x"73",x"87"),
  2073 => (x"c2",x"91",x"29",x"b7"),
  2074 => (x"73",x"81",x"ec",x"c2"),
  2075 => (x"c2",x"9a",x"cf",x"4a"),
  2076 => (x"72",x"48",x"c3",x"92"),
  2077 => (x"48",x"4a",x"70",x"30"),
  2078 => (x"79",x"70",x"b0",x"69"),
  2079 => (x"48",x"e8",x"c2",x"c2"),
  2080 => (x"c2",x"c2",x"78",x"c0"),
  2081 => (x"78",x"c0",x"48",x"e4"),
  2082 => (x"49",x"ea",x"fe",x"c2"),
  2083 => (x"70",x"87",x"cf",x"fa"),
  2084 => (x"aa",x"b7",x"c0",x"4a"),
  2085 => (x"87",x"f4",x"fd",x"03"),
  2086 => (x"87",x"c4",x"48",x"c0"),
  2087 => (x"4c",x"26",x"4d",x"26"),
  2088 => (x"4f",x"26",x"4b",x"26"),
  2089 => (x"00",x"00",x"00",x"00"),
  2090 => (x"00",x"00",x"00",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"00",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"00",x"00"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"00",x"00",x"00",x"00"),
  2096 => (x"00",x"00",x"00",x"00"),
  2097 => (x"00",x"00",x"00",x"00"),
  2098 => (x"00",x"00",x"00",x"00"),
  2099 => (x"00",x"00",x"00",x"00"),
  2100 => (x"00",x"00",x"00",x"00"),
  2101 => (x"00",x"00",x"00",x"00"),
  2102 => (x"00",x"00",x"00",x"00"),
  2103 => (x"00",x"00",x"00",x"00"),
  2104 => (x"00",x"00",x"00",x"00"),
  2105 => (x"00",x"00",x"00",x"00"),
  2106 => (x"00",x"00",x"00",x"00"),
  2107 => (x"72",x"4a",x"c0",x"1e"),
  2108 => (x"c2",x"91",x"c4",x"49"),
  2109 => (x"c0",x"81",x"ec",x"c2"),
  2110 => (x"d0",x"82",x"c1",x"79"),
  2111 => (x"ee",x"04",x"aa",x"b7"),
  2112 => (x"0e",x"4f",x"26",x"87"),
  2113 => (x"5d",x"5c",x"5b",x"5e"),
  2114 => (x"f6",x"4d",x"71",x"0e"),
  2115 => (x"4a",x"75",x"87",x"cb"),
  2116 => (x"92",x"2a",x"b7",x"c4"),
  2117 => (x"82",x"ec",x"c2",x"c2"),
  2118 => (x"9c",x"cf",x"4c",x"75"),
  2119 => (x"49",x"6a",x"94",x"c2"),
  2120 => (x"c3",x"2b",x"74",x"4b"),
  2121 => (x"74",x"48",x"c2",x"9b"),
  2122 => (x"ff",x"4c",x"70",x"30"),
  2123 => (x"71",x"48",x"74",x"bc"),
  2124 => (x"f5",x"7a",x"70",x"98"),
  2125 => (x"48",x"73",x"87",x"db"),
  2126 => (x"1e",x"87",x"e1",x"fd"),
  2127 => (x"bf",x"d0",x"ff",x"1e"),
  2128 => (x"c0",x"c0",x"c8",x"48"),
  2129 => (x"58",x"a6",x"c4",x"98"),
  2130 => (x"d0",x"02",x"98",x"70"),
  2131 => (x"bf",x"d0",x"ff",x"87"),
  2132 => (x"c0",x"c0",x"c8",x"48"),
  2133 => (x"58",x"a6",x"c4",x"98"),
  2134 => (x"f0",x"05",x"98",x"70"),
  2135 => (x"48",x"d0",x"ff",x"87"),
  2136 => (x"71",x"78",x"e1",x"c4"),
  2137 => (x"08",x"d4",x"ff",x"48"),
  2138 => (x"48",x"66",x"c8",x"78"),
  2139 => (x"78",x"08",x"d4",x"ff"),
  2140 => (x"1e",x"4f",x"26",x"26"),
  2141 => (x"c8",x"4a",x"71",x"1e"),
  2142 => (x"72",x"1e",x"49",x"66"),
  2143 => (x"87",x"fb",x"fe",x"49"),
  2144 => (x"d0",x"ff",x"86",x"c4"),
  2145 => (x"c0",x"c8",x"48",x"bf"),
  2146 => (x"a6",x"c4",x"98",x"c0"),
  2147 => (x"02",x"98",x"70",x"58"),
  2148 => (x"d0",x"ff",x"87",x"d0"),
  2149 => (x"c0",x"c8",x"48",x"bf"),
  2150 => (x"a6",x"c4",x"98",x"c0"),
  2151 => (x"05",x"98",x"70",x"58"),
  2152 => (x"d0",x"ff",x"87",x"f0"),
  2153 => (x"78",x"e0",x"c0",x"48"),
  2154 => (x"1e",x"4f",x"26",x"26"),
  2155 => (x"4b",x"71",x"1e",x"73"),
  2156 => (x"73",x"1e",x"66",x"c8"),
  2157 => (x"a2",x"e0",x"c1",x"4a"),
  2158 => (x"87",x"f7",x"fe",x"49"),
  2159 => (x"26",x"87",x"c4",x"26"),
  2160 => (x"26",x"4c",x"26",x"4d"),
  2161 => (x"1e",x"4f",x"26",x"4b"),
  2162 => (x"bf",x"d0",x"ff",x"1e"),
  2163 => (x"c0",x"c0",x"c8",x"48"),
  2164 => (x"58",x"a6",x"c4",x"98"),
  2165 => (x"d0",x"02",x"98",x"70"),
  2166 => (x"bf",x"d0",x"ff",x"87"),
  2167 => (x"c0",x"c0",x"c8",x"48"),
  2168 => (x"58",x"a6",x"c4",x"98"),
  2169 => (x"f0",x"05",x"98",x"70"),
  2170 => (x"48",x"d0",x"ff",x"87"),
  2171 => (x"71",x"78",x"c9",x"c4"),
  2172 => (x"08",x"d4",x"ff",x"48"),
  2173 => (x"4f",x"26",x"26",x"78"),
  2174 => (x"4a",x"71",x"1e",x"1e"),
  2175 => (x"87",x"c7",x"ff",x"49"),
  2176 => (x"48",x"bf",x"d0",x"ff"),
  2177 => (x"98",x"c0",x"c0",x"c8"),
  2178 => (x"70",x"58",x"a6",x"c4"),
  2179 => (x"87",x"d0",x"02",x"98"),
  2180 => (x"48",x"bf",x"d0",x"ff"),
  2181 => (x"98",x"c0",x"c0",x"c8"),
  2182 => (x"70",x"58",x"a6",x"c4"),
  2183 => (x"87",x"f0",x"05",x"98"),
  2184 => (x"c8",x"48",x"d0",x"ff"),
  2185 => (x"4f",x"26",x"26",x"78"),
  2186 => (x"1e",x"1e",x"73",x"1e"),
  2187 => (x"c1",x"c3",x"4b",x"71"),
  2188 => (x"c3",x"02",x"bf",x"c6"),
  2189 => (x"87",x"cc",x"c3",x"87"),
  2190 => (x"48",x"bf",x"d0",x"ff"),
  2191 => (x"98",x"c0",x"c0",x"c8"),
  2192 => (x"70",x"58",x"a6",x"c4"),
  2193 => (x"87",x"d0",x"02",x"98"),
  2194 => (x"48",x"bf",x"d0",x"ff"),
  2195 => (x"98",x"c0",x"c0",x"c8"),
  2196 => (x"70",x"58",x"a6",x"c4"),
  2197 => (x"87",x"f0",x"05",x"98"),
  2198 => (x"c4",x"48",x"d0",x"ff"),
  2199 => (x"48",x"73",x"78",x"c9"),
  2200 => (x"ff",x"b0",x"e0",x"c0"),
  2201 => (x"c3",x"78",x"08",x"d4"),
  2202 => (x"c0",x"48",x"fa",x"c0"),
  2203 => (x"02",x"66",x"cc",x"78"),
  2204 => (x"ff",x"c3",x"87",x"c5"),
  2205 => (x"c0",x"87",x"c2",x"49"),
  2206 => (x"c2",x"c1",x"c3",x"49"),
  2207 => (x"02",x"66",x"d0",x"59"),
  2208 => (x"d5",x"c5",x"87",x"c6"),
  2209 => (x"87",x"c4",x"4a",x"d5"),
  2210 => (x"4a",x"ff",x"ff",x"cf"),
  2211 => (x"5a",x"c6",x"c1",x"c3"),
  2212 => (x"48",x"c6",x"c1",x"c3"),
  2213 => (x"c4",x"26",x"78",x"c1"),
  2214 => (x"26",x"4d",x"26",x"87"),
  2215 => (x"26",x"4b",x"26",x"4c"),
  2216 => (x"5b",x"5e",x"0e",x"4f"),
  2217 => (x"71",x"0e",x"5d",x"5c"),
  2218 => (x"c2",x"c1",x"c3",x"4a"),
  2219 => (x"9a",x"72",x"4c",x"bf"),
  2220 => (x"49",x"87",x"cb",x"02"),
  2221 => (x"c9",x"c2",x"91",x"c8"),
  2222 => (x"83",x"71",x"4b",x"e2"),
  2223 => (x"cd",x"c2",x"87",x"c4"),
  2224 => (x"4d",x"c0",x"4b",x"e2"),
  2225 => (x"99",x"74",x"49",x"13"),
  2226 => (x"bf",x"fe",x"c0",x"c3"),
  2227 => (x"ff",x"b8",x"71",x"48"),
  2228 => (x"c1",x"78",x"08",x"d4"),
  2229 => (x"c8",x"85",x"2c",x"b7"),
  2230 => (x"e7",x"04",x"ad",x"b7"),
  2231 => (x"fa",x"c0",x"c3",x"87"),
  2232 => (x"80",x"c8",x"48",x"bf"),
  2233 => (x"58",x"fe",x"c0",x"c3"),
  2234 => (x"1e",x"87",x"ee",x"fe"),
  2235 => (x"4b",x"71",x"1e",x"73"),
  2236 => (x"02",x"9a",x"4a",x"13"),
  2237 => (x"49",x"72",x"87",x"cb"),
  2238 => (x"13",x"87",x"e6",x"fe"),
  2239 => (x"f5",x"05",x"9a",x"4a"),
  2240 => (x"87",x"d9",x"fe",x"87"),
  2241 => (x"c0",x"c3",x"1e",x"1e"),
  2242 => (x"c3",x"49",x"bf",x"fa"),
  2243 => (x"c1",x"48",x"fa",x"c0"),
  2244 => (x"c0",x"c4",x"78",x"a1"),
  2245 => (x"db",x"03",x"a9",x"b7"),
  2246 => (x"48",x"d4",x"ff",x"87"),
  2247 => (x"bf",x"fe",x"c0",x"c3"),
  2248 => (x"fa",x"c0",x"c3",x"78"),
  2249 => (x"c0",x"c3",x"49",x"bf"),
  2250 => (x"a1",x"c1",x"48",x"fa"),
  2251 => (x"b7",x"c0",x"c4",x"78"),
  2252 => (x"87",x"e5",x"04",x"a9"),
  2253 => (x"48",x"bf",x"d0",x"ff"),
  2254 => (x"98",x"c0",x"c0",x"c8"),
  2255 => (x"70",x"58",x"a6",x"c4"),
  2256 => (x"87",x"d0",x"02",x"98"),
  2257 => (x"48",x"bf",x"d0",x"ff"),
  2258 => (x"98",x"c0",x"c0",x"c8"),
  2259 => (x"70",x"58",x"a6",x"c4"),
  2260 => (x"87",x"f0",x"05",x"98"),
  2261 => (x"c8",x"48",x"d0",x"ff"),
  2262 => (x"c6",x"c1",x"c3",x"78"),
  2263 => (x"26",x"78",x"c0",x"48"),
  2264 => (x"00",x"00",x"4f",x"26"),
  2265 => (x"00",x"00",x"00",x"00"),
  2266 => (x"00",x"00",x"00",x"00"),
  2267 => (x"00",x"5f",x"5f",x"00"),
  2268 => (x"03",x"00",x"00",x"00"),
  2269 => (x"03",x"03",x"00",x"03"),
  2270 => (x"7f",x"14",x"00",x"00"),
  2271 => (x"7f",x"7f",x"14",x"7f"),
  2272 => (x"24",x"00",x"00",x"14"),
  2273 => (x"3a",x"6b",x"6b",x"2e"),
  2274 => (x"6a",x"4c",x"00",x"12"),
  2275 => (x"56",x"6c",x"18",x"36"),
  2276 => (x"7e",x"30",x"00",x"32"),
  2277 => (x"3a",x"77",x"59",x"4f"),
  2278 => (x"00",x"00",x"40",x"68"),
  2279 => (x"00",x"03",x"07",x"04"),
  2280 => (x"00",x"00",x"00",x"00"),
  2281 => (x"41",x"63",x"3e",x"1c"),
  2282 => (x"00",x"00",x"00",x"00"),
  2283 => (x"1c",x"3e",x"63",x"41"),
  2284 => (x"2a",x"08",x"00",x"00"),
  2285 => (x"3e",x"1c",x"1c",x"3e"),
  2286 => (x"08",x"00",x"08",x"2a"),
  2287 => (x"08",x"3e",x"3e",x"08"),
  2288 => (x"00",x"00",x"00",x"08"),
  2289 => (x"00",x"60",x"e0",x"80"),
  2290 => (x"08",x"00",x"00",x"00"),
  2291 => (x"08",x"08",x"08",x"08"),
  2292 => (x"00",x"00",x"00",x"08"),
  2293 => (x"00",x"60",x"60",x"00"),
  2294 => (x"60",x"40",x"00",x"00"),
  2295 => (x"06",x"0c",x"18",x"30"),
  2296 => (x"3e",x"00",x"01",x"03"),
  2297 => (x"7f",x"4d",x"59",x"7f"),
  2298 => (x"04",x"00",x"00",x"3e"),
  2299 => (x"00",x"7f",x"7f",x"06"),
  2300 => (x"42",x"00",x"00",x"00"),
  2301 => (x"4f",x"59",x"71",x"63"),
  2302 => (x"22",x"00",x"00",x"46"),
  2303 => (x"7f",x"49",x"49",x"63"),
  2304 => (x"1c",x"18",x"00",x"36"),
  2305 => (x"7f",x"7f",x"13",x"16"),
  2306 => (x"27",x"00",x"00",x"10"),
  2307 => (x"7d",x"45",x"45",x"67"),
  2308 => (x"3c",x"00",x"00",x"39"),
  2309 => (x"79",x"49",x"4b",x"7e"),
  2310 => (x"01",x"00",x"00",x"30"),
  2311 => (x"0f",x"79",x"71",x"01"),
  2312 => (x"36",x"00",x"00",x"07"),
  2313 => (x"7f",x"49",x"49",x"7f"),
  2314 => (x"06",x"00",x"00",x"36"),
  2315 => (x"3f",x"69",x"49",x"4f"),
  2316 => (x"00",x"00",x"00",x"1e"),
  2317 => (x"00",x"66",x"66",x"00"),
  2318 => (x"00",x"00",x"00",x"00"),
  2319 => (x"00",x"66",x"e6",x"80"),
  2320 => (x"08",x"00",x"00",x"00"),
  2321 => (x"22",x"14",x"14",x"08"),
  2322 => (x"14",x"00",x"00",x"22"),
  2323 => (x"14",x"14",x"14",x"14"),
  2324 => (x"22",x"00",x"00",x"14"),
  2325 => (x"08",x"14",x"14",x"22"),
  2326 => (x"02",x"00",x"00",x"08"),
  2327 => (x"0f",x"59",x"51",x"03"),
  2328 => (x"7f",x"3e",x"00",x"06"),
  2329 => (x"1f",x"55",x"5d",x"41"),
  2330 => (x"7e",x"00",x"00",x"1e"),
  2331 => (x"7f",x"09",x"09",x"7f"),
  2332 => (x"7f",x"00",x"00",x"7e"),
  2333 => (x"7f",x"49",x"49",x"7f"),
  2334 => (x"1c",x"00",x"00",x"36"),
  2335 => (x"41",x"41",x"63",x"3e"),
  2336 => (x"7f",x"00",x"00",x"41"),
  2337 => (x"3e",x"63",x"41",x"7f"),
  2338 => (x"7f",x"00",x"00",x"1c"),
  2339 => (x"41",x"49",x"49",x"7f"),
  2340 => (x"7f",x"00",x"00",x"41"),
  2341 => (x"01",x"09",x"09",x"7f"),
  2342 => (x"3e",x"00",x"00",x"01"),
  2343 => (x"7b",x"49",x"41",x"7f"),
  2344 => (x"7f",x"00",x"00",x"7a"),
  2345 => (x"7f",x"08",x"08",x"7f"),
  2346 => (x"00",x"00",x"00",x"7f"),
  2347 => (x"41",x"7f",x"7f",x"41"),
  2348 => (x"20",x"00",x"00",x"00"),
  2349 => (x"7f",x"40",x"40",x"60"),
  2350 => (x"7f",x"7f",x"00",x"3f"),
  2351 => (x"63",x"36",x"1c",x"08"),
  2352 => (x"7f",x"00",x"00",x"41"),
  2353 => (x"40",x"40",x"40",x"7f"),
  2354 => (x"7f",x"7f",x"00",x"40"),
  2355 => (x"7f",x"06",x"0c",x"06"),
  2356 => (x"7f",x"7f",x"00",x"7f"),
  2357 => (x"7f",x"18",x"0c",x"06"),
  2358 => (x"3e",x"00",x"00",x"7f"),
  2359 => (x"7f",x"41",x"41",x"7f"),
  2360 => (x"7f",x"00",x"00",x"3e"),
  2361 => (x"0f",x"09",x"09",x"7f"),
  2362 => (x"7f",x"3e",x"00",x"06"),
  2363 => (x"7e",x"7f",x"61",x"41"),
  2364 => (x"7f",x"00",x"00",x"40"),
  2365 => (x"7f",x"19",x"09",x"7f"),
  2366 => (x"26",x"00",x"00",x"66"),
  2367 => (x"7b",x"59",x"4d",x"6f"),
  2368 => (x"01",x"00",x"00",x"32"),
  2369 => (x"01",x"7f",x"7f",x"01"),
  2370 => (x"3f",x"00",x"00",x"01"),
  2371 => (x"7f",x"40",x"40",x"7f"),
  2372 => (x"0f",x"00",x"00",x"3f"),
  2373 => (x"3f",x"70",x"70",x"3f"),
  2374 => (x"7f",x"7f",x"00",x"0f"),
  2375 => (x"7f",x"30",x"18",x"30"),
  2376 => (x"63",x"41",x"00",x"7f"),
  2377 => (x"36",x"1c",x"1c",x"36"),
  2378 => (x"03",x"01",x"41",x"63"),
  2379 => (x"06",x"7c",x"7c",x"06"),
  2380 => (x"71",x"61",x"01",x"03"),
  2381 => (x"43",x"47",x"4d",x"59"),
  2382 => (x"00",x"00",x"00",x"41"),
  2383 => (x"41",x"41",x"7f",x"7f"),
  2384 => (x"03",x"01",x"00",x"00"),
  2385 => (x"30",x"18",x"0c",x"06"),
  2386 => (x"00",x"00",x"40",x"60"),
  2387 => (x"7f",x"7f",x"41",x"41"),
  2388 => (x"0c",x"08",x"00",x"00"),
  2389 => (x"0c",x"06",x"03",x"06"),
  2390 => (x"80",x"80",x"00",x"08"),
  2391 => (x"80",x"80",x"80",x"80"),
  2392 => (x"00",x"00",x"00",x"80"),
  2393 => (x"04",x"07",x"03",x"00"),
  2394 => (x"20",x"00",x"00",x"00"),
  2395 => (x"7c",x"54",x"54",x"74"),
  2396 => (x"7f",x"00",x"00",x"78"),
  2397 => (x"7c",x"44",x"44",x"7f"),
  2398 => (x"38",x"00",x"00",x"38"),
  2399 => (x"44",x"44",x"44",x"7c"),
  2400 => (x"38",x"00",x"00",x"00"),
  2401 => (x"7f",x"44",x"44",x"7c"),
  2402 => (x"38",x"00",x"00",x"7f"),
  2403 => (x"5c",x"54",x"54",x"7c"),
  2404 => (x"04",x"00",x"00",x"18"),
  2405 => (x"05",x"05",x"7f",x"7e"),
  2406 => (x"18",x"00",x"00",x"00"),
  2407 => (x"fc",x"a4",x"a4",x"bc"),
  2408 => (x"7f",x"00",x"00",x"7c"),
  2409 => (x"7c",x"04",x"04",x"7f"),
  2410 => (x"00",x"00",x"00",x"78"),
  2411 => (x"40",x"7d",x"3d",x"00"),
  2412 => (x"80",x"00",x"00",x"00"),
  2413 => (x"7d",x"fd",x"80",x"80"),
  2414 => (x"7f",x"00",x"00",x"00"),
  2415 => (x"6c",x"38",x"10",x"7f"),
  2416 => (x"00",x"00",x"00",x"44"),
  2417 => (x"40",x"7f",x"3f",x"00"),
  2418 => (x"7c",x"7c",x"00",x"00"),
  2419 => (x"7c",x"0c",x"18",x"0c"),
  2420 => (x"7c",x"00",x"00",x"78"),
  2421 => (x"7c",x"04",x"04",x"7c"),
  2422 => (x"38",x"00",x"00",x"78"),
  2423 => (x"7c",x"44",x"44",x"7c"),
  2424 => (x"fc",x"00",x"00",x"38"),
  2425 => (x"3c",x"24",x"24",x"fc"),
  2426 => (x"18",x"00",x"00",x"18"),
  2427 => (x"fc",x"24",x"24",x"3c"),
  2428 => (x"7c",x"00",x"00",x"fc"),
  2429 => (x"0c",x"04",x"04",x"7c"),
  2430 => (x"48",x"00",x"00",x"08"),
  2431 => (x"74",x"54",x"54",x"5c"),
  2432 => (x"04",x"00",x"00",x"20"),
  2433 => (x"44",x"44",x"7f",x"3f"),
  2434 => (x"3c",x"00",x"00",x"00"),
  2435 => (x"7c",x"40",x"40",x"7c"),
  2436 => (x"1c",x"00",x"00",x"7c"),
  2437 => (x"3c",x"60",x"60",x"3c"),
  2438 => (x"7c",x"3c",x"00",x"1c"),
  2439 => (x"7c",x"60",x"30",x"60"),
  2440 => (x"6c",x"44",x"00",x"3c"),
  2441 => (x"6c",x"38",x"10",x"38"),
  2442 => (x"1c",x"00",x"00",x"44"),
  2443 => (x"3c",x"60",x"e0",x"bc"),
  2444 => (x"44",x"00",x"00",x"1c"),
  2445 => (x"4c",x"5c",x"74",x"64"),
  2446 => (x"08",x"00",x"00",x"44"),
  2447 => (x"41",x"77",x"3e",x"08"),
  2448 => (x"00",x"00",x"00",x"41"),
  2449 => (x"00",x"7f",x"7f",x"00"),
  2450 => (x"41",x"00",x"00",x"00"),
  2451 => (x"08",x"3e",x"77",x"41"),
  2452 => (x"01",x"02",x"00",x"08"),
  2453 => (x"02",x"02",x"03",x"01"),
  2454 => (x"7f",x"7f",x"00",x"01"),
  2455 => (x"7f",x"7f",x"7f",x"7f"),
  2456 => (x"08",x"08",x"00",x"7f"),
  2457 => (x"3e",x"3e",x"1c",x"1c"),
  2458 => (x"7f",x"7f",x"7f",x"7f"),
  2459 => (x"1c",x"1c",x"3e",x"3e"),
  2460 => (x"10",x"00",x"08",x"08"),
  2461 => (x"18",x"7c",x"7c",x"18"),
  2462 => (x"10",x"00",x"00",x"10"),
  2463 => (x"30",x"7c",x"7c",x"30"),
  2464 => (x"30",x"10",x"00",x"10"),
  2465 => (x"1e",x"78",x"60",x"60"),
  2466 => (x"66",x"42",x"00",x"06"),
  2467 => (x"66",x"3c",x"18",x"3c"),
  2468 => (x"38",x"78",x"00",x"42"),
  2469 => (x"6c",x"c6",x"c2",x"6a"),
  2470 => (x"00",x"60",x"00",x"38"),
  2471 => (x"00",x"00",x"60",x"00"),
  2472 => (x"5e",x"0e",x"00",x"60"),
  2473 => (x"0e",x"5d",x"5c",x"5b"),
  2474 => (x"c3",x"4c",x"71",x"1e"),
  2475 => (x"4b",x"bf",x"ce",x"c1"),
  2476 => (x"48",x"d2",x"c1",x"c3"),
  2477 => (x"1e",x"74",x"78",x"c0"),
  2478 => (x"1e",x"fd",x"dc",x"c2"),
  2479 => (x"87",x"fc",x"e6",x"fd"),
  2480 => (x"6b",x"97",x"86",x"c8"),
  2481 => (x"c1",x"02",x"99",x"49"),
  2482 => (x"1e",x"c0",x"87",x"c6"),
  2483 => (x"c3",x"48",x"a6",x"c4"),
  2484 => (x"78",x"bf",x"d2",x"c1"),
  2485 => (x"02",x"ac",x"66",x"c4"),
  2486 => (x"4d",x"c0",x"87",x"c4"),
  2487 => (x"4d",x"c1",x"87",x"c2"),
  2488 => (x"66",x"c8",x"1e",x"75"),
  2489 => (x"87",x"c0",x"ed",x"49"),
  2490 => (x"e0",x"c0",x"86",x"c8"),
  2491 => (x"87",x"f1",x"ee",x"49"),
  2492 => (x"6a",x"4a",x"a3",x"c4"),
  2493 => (x"87",x"f3",x"ef",x"49"),
  2494 => (x"c3",x"87",x"c9",x"f0"),
  2495 => (x"48",x"bf",x"d2",x"c1"),
  2496 => (x"c1",x"c3",x"80",x"c1"),
  2497 => (x"83",x"cc",x"58",x"d6"),
  2498 => (x"99",x"49",x"6b",x"97"),
  2499 => (x"87",x"fa",x"fe",x"05"),
  2500 => (x"bf",x"d2",x"c1",x"c3"),
  2501 => (x"ad",x"b7",x"c8",x"4d"),
  2502 => (x"c0",x"87",x"d9",x"03"),
  2503 => (x"c1",x"c3",x"1e",x"1e"),
  2504 => (x"ec",x"49",x"bf",x"d2"),
  2505 => (x"86",x"c8",x"87",x"c2"),
  2506 => (x"c1",x"87",x"d9",x"ef"),
  2507 => (x"ad",x"b7",x"c8",x"85"),
  2508 => (x"87",x"e7",x"ff",x"04"),
  2509 => (x"26",x"4d",x"26",x"26"),
  2510 => (x"26",x"4b",x"26",x"4c"),
  2511 => (x"67",x"69",x"48",x"4f"),
  2512 => (x"67",x"69",x"6c",x"68"),
  2513 => (x"72",x"20",x"74",x"68"),
  2514 => (x"25",x"20",x"77",x"6f"),
  2515 => (x"4d",x"00",x"0a",x"64"),
  2516 => (x"20",x"75",x"6e",x"65"),
  2517 => (x"69",x"73",x"69",x"76"),
  2518 => (x"20",x"65",x"6c",x"62"),
  2519 => (x"00",x"0a",x"64",x"25"),
  2520 => (x"6c",x"6c",x"61",x"43"),
  2521 => (x"6b",x"63",x"61",x"62"),
  2522 => (x"0a",x"78",x"25",x"20"),
  2523 => (x"4a",x"71",x"1e",x"00"),
  2524 => (x"5a",x"d2",x"c1",x"c3"),
  2525 => (x"bf",x"d6",x"c1",x"c3"),
  2526 => (x"87",x"e6",x"fc",x"49"),
  2527 => (x"bf",x"d2",x"c1",x"c3"),
  2528 => (x"c3",x"89",x"c1",x"49"),
  2529 => (x"71",x"59",x"da",x"c1"),
  2530 => (x"26",x"87",x"d7",x"fc"),
  2531 => (x"c0",x"c1",x"1e",x"4f"),
  2532 => (x"87",x"e4",x"e9",x"49"),
  2533 => (x"48",x"c1",x"ec",x"c2"),
  2534 => (x"4f",x"26",x"78",x"c0"),
  2535 => (x"5c",x"5b",x"5e",x"0e"),
  2536 => (x"86",x"f4",x"0e",x"5d"),
  2537 => (x"c0",x"48",x"a6",x"c8"),
  2538 => (x"7e",x"bf",x"ec",x"78"),
  2539 => (x"c1",x"c3",x"80",x"fc"),
  2540 => (x"c3",x"78",x"bf",x"ce"),
  2541 => (x"4d",x"bf",x"da",x"c1"),
  2542 => (x"c7",x"4c",x"bf",x"e8"),
  2543 => (x"87",x"c3",x"e5",x"49"),
  2544 => (x"99",x"c2",x"49",x"70"),
  2545 => (x"c2",x"87",x"cf",x"05"),
  2546 => (x"49",x"bf",x"f9",x"eb"),
  2547 => (x"99",x"6e",x"b9",x"ff"),
  2548 => (x"c0",x"02",x"99",x"c1"),
  2549 => (x"49",x"c7",x"87",x"fd"),
  2550 => (x"70",x"87",x"e8",x"e4"),
  2551 => (x"87",x"cd",x"02",x"98"),
  2552 => (x"c7",x"87",x"d6",x"e0"),
  2553 => (x"87",x"db",x"e4",x"49"),
  2554 => (x"f3",x"05",x"98",x"70"),
  2555 => (x"c1",x"ec",x"c2",x"87"),
  2556 => (x"dd",x"c2",x"1e",x"bf"),
  2557 => (x"e2",x"fd",x"1e",x"cf"),
  2558 => (x"86",x"c8",x"87",x"c2"),
  2559 => (x"bf",x"c1",x"ec",x"c2"),
  2560 => (x"c2",x"ba",x"c1",x"4a"),
  2561 => (x"c1",x"5a",x"c5",x"ec"),
  2562 => (x"e7",x"49",x"a2",x"c0"),
  2563 => (x"a6",x"c8",x"87",x"ea"),
  2564 => (x"c2",x"78",x"c1",x"48"),
  2565 => (x"6e",x"48",x"f9",x"eb"),
  2566 => (x"c1",x"ec",x"c2",x"78"),
  2567 => (x"da",x"c1",x"05",x"bf"),
  2568 => (x"48",x"a6",x"c4",x"87"),
  2569 => (x"78",x"c0",x"c0",x"c8"),
  2570 => (x"7e",x"c5",x"ec",x"c2"),
  2571 => (x"49",x"bf",x"97",x"6e"),
  2572 => (x"80",x"c1",x"48",x"6e"),
  2573 => (x"71",x"58",x"a6",x"c4"),
  2574 => (x"70",x"87",x"c8",x"e3"),
  2575 => (x"87",x"c3",x"02",x"98"),
  2576 => (x"c4",x"b4",x"66",x"c4"),
  2577 => (x"b7",x"c1",x"48",x"66"),
  2578 => (x"58",x"a6",x"c8",x"28"),
  2579 => (x"ff",x"05",x"98",x"70"),
  2580 => (x"49",x"74",x"87",x"da"),
  2581 => (x"71",x"99",x"ff",x"c3"),
  2582 => (x"e5",x"49",x"c0",x"1e"),
  2583 => (x"49",x"74",x"87",x"cd"),
  2584 => (x"71",x"29",x"b7",x"c8"),
  2585 => (x"e5",x"49",x"c1",x"1e"),
  2586 => (x"86",x"c8",x"87",x"c1"),
  2587 => (x"e2",x"49",x"fd",x"c3"),
  2588 => (x"fa",x"c3",x"87",x"d1"),
  2589 => (x"87",x"cb",x"e2",x"49"),
  2590 => (x"74",x"87",x"e9",x"c9"),
  2591 => (x"99",x"ff",x"c3",x"49"),
  2592 => (x"71",x"2c",x"b7",x"c8"),
  2593 => (x"02",x"9c",x"74",x"b4"),
  2594 => (x"c8",x"ff",x"87",x"df"),
  2595 => (x"49",x"6e",x"7e",x"bf"),
  2596 => (x"bf",x"fd",x"eb",x"c2"),
  2597 => (x"a9",x"c0",x"c2",x"89"),
  2598 => (x"87",x"c4",x"c0",x"03"),
  2599 => (x"87",x"cf",x"4c",x"c0"),
  2600 => (x"48",x"fd",x"eb",x"c2"),
  2601 => (x"c6",x"c0",x"78",x"6e"),
  2602 => (x"fd",x"eb",x"c2",x"87"),
  2603 => (x"74",x"78",x"c0",x"48"),
  2604 => (x"05",x"99",x"c8",x"49"),
  2605 => (x"f5",x"c3",x"87",x"ce"),
  2606 => (x"87",x"c7",x"e1",x"49"),
  2607 => (x"99",x"c2",x"49",x"70"),
  2608 => (x"87",x"ee",x"c0",x"02"),
  2609 => (x"bf",x"d6",x"c1",x"c3"),
  2610 => (x"87",x"c9",x"c0",x"02"),
  2611 => (x"c3",x"88",x"c1",x"48"),
  2612 => (x"d8",x"58",x"da",x"c1"),
  2613 => (x"d2",x"c1",x"c3",x"87"),
  2614 => (x"91",x"cc",x"49",x"bf"),
  2615 => (x"c8",x"81",x"66",x"c4"),
  2616 => (x"bf",x"6e",x"7e",x"a1"),
  2617 => (x"87",x"c5",x"c0",x"02"),
  2618 => (x"73",x"49",x"ff",x"4b"),
  2619 => (x"48",x"a6",x"c8",x"0f"),
  2620 => (x"49",x"74",x"78",x"c1"),
  2621 => (x"c0",x"05",x"99",x"c4"),
  2622 => (x"f2",x"c3",x"87",x"ce"),
  2623 => (x"87",x"c3",x"e0",x"49"),
  2624 => (x"99",x"c2",x"49",x"70"),
  2625 => (x"87",x"fe",x"c0",x"02"),
  2626 => (x"c3",x"48",x"a6",x"c8"),
  2627 => (x"78",x"bf",x"d2",x"c1"),
  2628 => (x"c1",x"49",x"66",x"c8"),
  2629 => (x"d6",x"c1",x"c3",x"89"),
  2630 => (x"b7",x"6e",x"7e",x"bf"),
  2631 => (x"ca",x"c0",x"06",x"a9"),
  2632 => (x"80",x"c1",x"48",x"87"),
  2633 => (x"58",x"da",x"c1",x"c3"),
  2634 => (x"c8",x"87",x"d6",x"c0"),
  2635 => (x"91",x"cc",x"49",x"66"),
  2636 => (x"c8",x"81",x"66",x"c4"),
  2637 => (x"bf",x"6e",x"7e",x"a1"),
  2638 => (x"87",x"c5",x"c0",x"02"),
  2639 => (x"73",x"49",x"fe",x"4b"),
  2640 => (x"48",x"a6",x"c8",x"0f"),
  2641 => (x"fd",x"c3",x"78",x"c1"),
  2642 => (x"f6",x"de",x"ff",x"49"),
  2643 => (x"c2",x"49",x"70",x"87"),
  2644 => (x"ee",x"c0",x"02",x"99"),
  2645 => (x"d6",x"c1",x"c3",x"87"),
  2646 => (x"c9",x"c0",x"02",x"bf"),
  2647 => (x"d6",x"c1",x"c3",x"87"),
  2648 => (x"c0",x"78",x"c0",x"48"),
  2649 => (x"c1",x"c3",x"87",x"d8"),
  2650 => (x"cc",x"49",x"bf",x"d2"),
  2651 => (x"81",x"66",x"c4",x"91"),
  2652 => (x"6e",x"7e",x"a1",x"c8"),
  2653 => (x"c5",x"c0",x"02",x"bf"),
  2654 => (x"49",x"fd",x"4b",x"87"),
  2655 => (x"a6",x"c8",x"0f",x"73"),
  2656 => (x"c3",x"78",x"c1",x"48"),
  2657 => (x"dd",x"ff",x"49",x"fa"),
  2658 => (x"49",x"70",x"87",x"f9"),
  2659 => (x"c1",x"02",x"99",x"c2"),
  2660 => (x"a6",x"c8",x"87",x"c0"),
  2661 => (x"d2",x"c1",x"c3",x"48"),
  2662 => (x"66",x"c8",x"78",x"bf"),
  2663 => (x"c4",x"88",x"c1",x"48"),
  2664 => (x"c1",x"c3",x"58",x"a6"),
  2665 => (x"6e",x"48",x"bf",x"d6"),
  2666 => (x"c0",x"03",x"a8",x"b7"),
  2667 => (x"c1",x"c3",x"87",x"c9"),
  2668 => (x"78",x"6e",x"48",x"d6"),
  2669 => (x"c8",x"87",x"d6",x"c0"),
  2670 => (x"91",x"cc",x"49",x"66"),
  2671 => (x"c8",x"81",x"66",x"c4"),
  2672 => (x"bf",x"6e",x"7e",x"a1"),
  2673 => (x"87",x"c5",x"c0",x"02"),
  2674 => (x"73",x"49",x"fc",x"4b"),
  2675 => (x"48",x"a6",x"c8",x"0f"),
  2676 => (x"c1",x"c3",x"78",x"c1"),
  2677 => (x"c0",x"4b",x"bf",x"d6"),
  2678 => (x"c0",x"06",x"ab",x"b7"),
  2679 => (x"8b",x"c1",x"87",x"c9"),
  2680 => (x"01",x"ab",x"b7",x"c0"),
  2681 => (x"74",x"87",x"f7",x"ff"),
  2682 => (x"99",x"f0",x"c3",x"49"),
  2683 => (x"87",x"cf",x"c0",x"05"),
  2684 => (x"ff",x"49",x"da",x"c1"),
  2685 => (x"70",x"87",x"cc",x"dc"),
  2686 => (x"02",x"99",x"c2",x"49"),
  2687 => (x"c3",x"87",x"e8",x"c2"),
  2688 => (x"7e",x"bf",x"ce",x"c1"),
  2689 => (x"bf",x"d6",x"c1",x"c3"),
  2690 => (x"ab",x"b7",x"c0",x"4b"),
  2691 => (x"87",x"d0",x"c0",x"06"),
  2692 => (x"80",x"cc",x"48",x"6e"),
  2693 => (x"c1",x"58",x"a6",x"c4"),
  2694 => (x"ab",x"b7",x"c0",x"8b"),
  2695 => (x"87",x"f0",x"ff",x"01"),
  2696 => (x"4a",x"bf",x"97",x"6e"),
  2697 => (x"c0",x"02",x"8a",x"c1"),
  2698 => (x"02",x"8a",x"87",x"f7"),
  2699 => (x"8a",x"87",x"d6",x"c0"),
  2700 => (x"87",x"ca",x"c1",x"02"),
  2701 => (x"ee",x"c1",x"05",x"8a"),
  2702 => (x"c8",x"4a",x"6e",x"87"),
  2703 => (x"f4",x"49",x"6a",x"82"),
  2704 => (x"e2",x"c1",x"87",x"eb"),
  2705 => (x"c8",x"4b",x"6e",x"87"),
  2706 => (x"c2",x"1e",x"6b",x"83"),
  2707 => (x"fd",x"1e",x"e0",x"dd"),
  2708 => (x"c8",x"87",x"e9",x"d8"),
  2709 => (x"c3",x"4b",x"6b",x"86"),
  2710 => (x"49",x"bf",x"d6",x"c1"),
  2711 => (x"c6",x"c1",x"0f",x"73"),
  2712 => (x"c8",x"49",x"6e",x"87"),
  2713 => (x"69",x"48",x"c1",x"81"),
  2714 => (x"c3",x"49",x"70",x"30"),
  2715 => (x"48",x"bf",x"ca",x"c1"),
  2716 => (x"c1",x"c3",x"b8",x"71"),
  2717 => (x"a6",x"c8",x"58",x"ce"),
  2718 => (x"c0",x"78",x"c1",x"48"),
  2719 => (x"49",x"6e",x"87",x"e9"),
  2720 => (x"48",x"6e",x"81",x"c8"),
  2721 => (x"a6",x"c8",x"80",x"cb"),
  2722 => (x"97",x"66",x"c4",x"58"),
  2723 => (x"a2",x"c1",x"4a",x"bf"),
  2724 => (x"49",x"69",x"97",x"4b"),
  2725 => (x"c0",x"04",x"ab",x"b7"),
  2726 => (x"4b",x"c0",x"87",x"c2"),
  2727 => (x"97",x"0b",x"66",x"c4"),
  2728 => (x"a6",x"c8",x"0b",x"7b"),
  2729 => (x"75",x"78",x"c1",x"48"),
  2730 => (x"e9",x"c0",x"02",x"9d"),
  2731 => (x"c0",x"02",x"6d",x"87"),
  2732 => (x"49",x"6d",x"87",x"e4"),
  2733 => (x"87",x"cb",x"d9",x"ff"),
  2734 => (x"99",x"c1",x"49",x"70"),
  2735 => (x"87",x"cb",x"c0",x"02"),
  2736 => (x"c3",x"4b",x"a5",x"c4"),
  2737 => (x"49",x"bf",x"d6",x"c1"),
  2738 => (x"c8",x"0f",x"4b",x"6b"),
  2739 => (x"c5",x"c0",x"02",x"85"),
  2740 => (x"ff",x"05",x"6d",x"87"),
  2741 => (x"66",x"c8",x"87",x"dc"),
  2742 => (x"87",x"c8",x"c0",x"02"),
  2743 => (x"bf",x"d6",x"c1",x"c3"),
  2744 => (x"87",x"fe",x"ee",x"49"),
  2745 => (x"cc",x"f1",x"8e",x"f4"),
  2746 => (x"11",x"12",x"58",x"87"),
  2747 => (x"1c",x"1b",x"1d",x"14"),
  2748 => (x"91",x"59",x"5a",x"23"),
  2749 => (x"eb",x"f2",x"f5",x"94"),
  2750 => (x"00",x"00",x"00",x"f4"),
  2751 => (x"00",x"00",x"00",x"00"),
  2752 => (x"00",x"00",x"00",x"00"),
  2753 => (x"14",x"12",x"58",x"00"),
  2754 => (x"1c",x"1b",x"1d",x"11"),
  2755 => (x"94",x"59",x"5a",x"23"),
  2756 => (x"eb",x"f2",x"f5",x"91"),
  2757 => (x"00",x"00",x"00",x"f4"),
  2758 => (x"00",x"00",x"2b",x"1c"),
  2759 => (x"4f",x"54",x"55",x"41"),
  2760 => (x"54",x"4f",x"4f",x"42"),
  2761 => (x"00",x"53",x"45",x"4e"),
  2762 => (x"00",x"00",x"1e",x"78"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

